magic
tech sky130A
magscale 1 2
timestamp 1655578206
<< metal1 >>
rect 3878 700748 3884 700800
rect 3936 700788 3942 700800
rect 8110 700788 8116 700800
rect 3936 700760 8116 700788
rect 3936 700748 3942 700760
rect 8110 700748 8116 700760
rect 8168 700748 8174 700800
rect 348786 700544 348792 700596
rect 348844 700584 348850 700596
rect 355870 700584 355876 700596
rect 348844 700556 355876 700584
rect 348844 700544 348850 700556
rect 355870 700544 355876 700556
rect 355928 700544 355934 700596
rect 105446 700272 105452 700324
rect 105504 700312 105510 700324
rect 113910 700312 113916 700324
rect 105504 700284 113916 700312
rect 105504 700272 105510 700284
rect 113910 700272 113916 700284
rect 113968 700272 113974 700324
rect 170306 700272 170312 700324
rect 170364 700312 170370 700324
rect 179874 700312 179880 700324
rect 170364 700284 179880 700312
rect 170364 700272 170370 700284
rect 179874 700272 179880 700284
rect 179932 700272 179938 700324
rect 218974 700272 218980 700324
rect 219032 700312 219038 700324
rect 223850 700312 223856 700324
rect 219032 700284 223856 700312
rect 219032 700272 219038 700284
rect 223850 700272 223856 700284
rect 223908 700272 223914 700324
rect 235166 700272 235172 700324
rect 235224 700312 235230 700324
rect 245838 700312 245844 700324
rect 235224 700284 245844 700312
rect 235224 700272 235230 700284
rect 245838 700272 245844 700284
rect 245896 700272 245902 700324
rect 283834 700272 283840 700324
rect 283892 700312 283898 700324
rect 289814 700312 289820 700324
rect 283892 700284 289820 700312
rect 283892 700272 283898 700284
rect 289814 700272 289820 700284
rect 289872 700272 289878 700324
rect 300118 700272 300124 700324
rect 300176 700312 300182 700324
rect 311894 700312 311900 700324
rect 300176 700284 311900 700312
rect 300176 700272 300182 700284
rect 311894 700272 311900 700284
rect 311952 700272 311958 700324
rect 364978 700272 364984 700324
rect 365036 700312 365042 700324
rect 377858 700312 377864 700324
rect 365036 700284 377864 700312
rect 365036 700272 365042 700284
rect 377858 700272 377864 700284
rect 377916 700272 377922 700324
rect 429838 700272 429844 700324
rect 429896 700312 429902 700324
rect 443822 700312 443828 700324
rect 429896 700284 443828 700312
rect 429896 700272 429902 700284
rect 443822 700272 443828 700284
rect 443880 700272 443886 700324
rect 478506 700272 478512 700324
rect 478564 700312 478570 700324
rect 487798 700312 487804 700324
rect 478564 700284 487804 700312
rect 478564 700272 478570 700284
rect 487798 700272 487804 700284
rect 487856 700272 487862 700324
rect 494790 700272 494796 700324
rect 494848 700312 494854 700324
rect 509786 700312 509792 700324
rect 494848 700284 509792 700312
rect 494848 700272 494854 700284
rect 509786 700272 509792 700284
rect 509844 700272 509850 700324
rect 527174 700272 527180 700324
rect 527232 700312 527238 700324
rect 531774 700312 531780 700324
rect 527232 700284 531780 700312
rect 527232 700272 527238 700284
rect 531774 700272 531780 700284
rect 531832 700272 531838 700324
rect 543458 700272 543464 700324
rect 543516 700312 543522 700324
rect 553762 700312 553768 700324
rect 543516 700284 553768 700312
rect 543516 700272 543522 700284
rect 553762 700272 553768 700284
rect 553820 700272 553826 700324
rect 559650 700272 559656 700324
rect 559708 700312 559714 700324
rect 575750 700312 575756 700324
rect 559708 700284 575756 700312
rect 559708 700272 559714 700284
rect 575750 700272 575756 700284
rect 575808 700272 575814 700324
rect 24302 700204 24308 700256
rect 24360 700244 24366 700256
rect 25958 700244 25964 700256
rect 24360 700216 25964 700244
rect 24360 700204 24366 700216
rect 25958 700204 25964 700216
rect 26016 700204 26022 700256
rect 40494 700204 40500 700256
rect 40552 700244 40558 700256
rect 47946 700244 47952 700256
rect 40552 700216 47952 700244
rect 40552 700204 40558 700216
rect 47946 700204 47952 700216
rect 48004 700204 48010 700256
rect 70026 700204 70032 700256
rect 70084 700244 70090 700256
rect 72970 700244 72976 700256
rect 70084 700216 72976 700244
rect 70084 700204 70090 700216
rect 72970 700204 72976 700216
rect 73028 700204 73034 700256
rect 89162 700204 89168 700256
rect 89220 700244 89226 700256
rect 91922 700244 91928 700256
rect 89220 700216 91928 700244
rect 89220 700204 89226 700216
rect 91922 700204 91928 700216
rect 91980 700204 91986 700256
rect 135990 700204 135996 700256
rect 136048 700244 136054 700256
rect 137830 700244 137836 700256
rect 136048 700216 137836 700244
rect 136048 700204 136054 700216
rect 137830 700204 137836 700216
rect 137888 700204 137894 700256
rect 154114 700204 154120 700256
rect 154172 700244 154178 700256
rect 157886 700244 157892 700256
rect 154172 700216 157892 700244
rect 154172 700204 154178 700216
rect 157886 700204 157892 700216
rect 157944 700204 157950 700256
rect 201954 700204 201960 700256
rect 202012 700244 202018 700256
rect 202782 700244 202788 700256
rect 202012 700216 202788 700244
rect 202012 700204 202018 700216
rect 202782 700204 202788 700216
rect 202840 700204 202846 700256
rect 397454 700204 397460 700256
rect 397512 700244 397518 700256
rect 399846 700244 399852 700256
rect 397512 700216 399852 700244
rect 397512 700204 397518 700216
rect 399846 700204 399852 700216
rect 399904 700204 399910 700256
rect 413646 700204 413652 700256
rect 413704 700244 413710 700256
rect 421834 700244 421840 700256
rect 413704 700216 421840 700244
rect 413704 700204 413710 700216
rect 421834 700204 421840 700216
rect 421892 700204 421898 700256
rect 462314 700204 462320 700256
rect 462372 700244 462378 700256
rect 465810 700244 465816 700256
rect 462372 700216 465816 700244
rect 462372 700204 462378 700216
rect 465810 700204 465816 700216
rect 465868 700204 465874 700256
rect 332502 700068 332508 700120
rect 332560 700108 332566 700120
rect 333882 700108 333888 700120
rect 332560 700080 333888 700108
rect 332560 700068 332566 700080
rect 333882 700068 333888 700080
rect 333940 700068 333946 700120
rect 578418 682456 578424 682508
rect 578476 682496 578482 682508
rect 579982 682496 579988 682508
rect 578476 682468 579988 682496
rect 578476 682456 578482 682468
rect 579982 682456 579988 682468
rect 580040 682456 580046 682508
rect 14 423580 20 423632
rect 72 423620 78 423632
rect 566 423620 572 423632
rect 72 423592 572 423620
rect 72 423580 78 423592
rect 566 423580 572 423592
rect 624 423580 630 423632
rect 578234 397468 578240 397520
rect 578292 397508 578298 397520
rect 580258 397508 580264 397520
rect 578292 397480 580264 397508
rect 578292 397468 578298 397480
rect 580258 397468 580264 397480
rect 580316 397468 580322 397520
rect 578326 351024 578332 351076
rect 578384 351064 578390 351076
rect 580258 351064 580264 351076
rect 578384 351036 580264 351064
rect 578384 351024 578390 351036
rect 580258 351024 580264 351036
rect 580316 351024 580322 351076
rect 578510 303696 578516 303748
rect 578568 303736 578574 303748
rect 580258 303736 580264 303748
rect 578568 303708 580264 303736
rect 578568 303696 578574 303708
rect 580258 303696 580264 303708
rect 580316 303696 580322 303748
rect 578878 273164 578884 273216
rect 578936 273204 578942 273216
rect 580810 273204 580816 273216
rect 578936 273176 580816 273204
rect 578936 273164 578942 273176
rect 580810 273164 580816 273176
rect 580868 273164 580874 273216
rect 578602 255280 578608 255332
rect 578660 255320 578666 255332
rect 580258 255320 580264 255332
rect 578660 255292 580264 255320
rect 578660 255280 578666 255292
rect 580258 255280 580264 255292
rect 580316 255280 580322 255332
rect 578326 208360 578332 208412
rect 578384 208400 578390 208412
rect 580258 208400 580264 208412
rect 578384 208372 580264 208400
rect 578384 208360 578390 208372
rect 580258 208360 580264 208372
rect 580316 208360 580322 208412
rect 578234 60664 578240 60716
rect 578292 60704 578298 60716
rect 580810 60704 580816 60716
rect 578292 60676 580816 60704
rect 578292 60664 578298 60676
rect 580810 60664 580816 60676
rect 580868 60664 580874 60716
rect 11146 3884 11152 3936
rect 11204 3924 11210 3936
rect 14502 3924 14508 3936
rect 11204 3896 14508 3924
rect 11204 3884 11210 3896
rect 14502 3884 14508 3896
rect 14560 3884 14566 3936
rect 14734 3884 14740 3936
rect 14792 3924 14798 3936
rect 17998 3924 18004 3936
rect 14792 3896 18004 3924
rect 14792 3884 14798 3896
rect 17998 3884 18004 3896
rect 18056 3884 18062 3936
rect 20622 3884 20628 3936
rect 20680 3924 20686 3936
rect 23794 3924 23800 3936
rect 20680 3896 23800 3924
rect 20680 3884 20686 3896
rect 23794 3884 23800 3896
rect 23852 3884 23858 3936
rect 24210 3884 24216 3936
rect 24268 3924 24274 3936
rect 27290 3924 27296 3936
rect 24268 3896 27296 3924
rect 24268 3884 24274 3896
rect 27290 3884 27296 3896
rect 27348 3884 27354 3936
rect 27706 3884 27712 3936
rect 27764 3924 27770 3936
rect 30694 3924 30700 3936
rect 27764 3896 30700 3924
rect 27764 3884 27770 3896
rect 30694 3884 30700 3896
rect 30752 3884 30758 3936
rect 32398 3884 32404 3936
rect 32456 3924 32462 3936
rect 35386 3924 35392 3936
rect 32456 3896 35392 3924
rect 32456 3884 32462 3896
rect 35386 3884 35392 3896
rect 35444 3884 35450 3936
rect 38378 3884 38384 3936
rect 38436 3924 38442 3936
rect 41182 3924 41188 3936
rect 38436 3896 41188 3924
rect 38436 3884 38442 3896
rect 41182 3884 41188 3896
rect 41240 3884 41246 3936
rect 43070 3884 43076 3936
rect 43128 3924 43134 3936
rect 45782 3924 45788 3936
rect 43128 3896 45788 3924
rect 43128 3884 43134 3896
rect 45782 3884 45788 3896
rect 45840 3884 45846 3936
rect 46658 3884 46664 3936
rect 46716 3924 46722 3936
rect 49278 3924 49284 3936
rect 46716 3896 49284 3924
rect 46716 3884 46722 3896
rect 49278 3884 49284 3896
rect 49336 3884 49342 3936
rect 50154 3884 50160 3936
rect 50212 3924 50218 3936
rect 52774 3924 52780 3936
rect 50212 3896 52780 3924
rect 50212 3884 50218 3896
rect 52774 3884 52780 3896
rect 52832 3884 52838 3936
rect 56042 3884 56048 3936
rect 56100 3924 56106 3936
rect 58570 3924 58576 3936
rect 56100 3896 58576 3924
rect 56100 3884 56106 3896
rect 58570 3884 58576 3896
rect 58628 3884 58634 3936
rect 72602 3884 72608 3936
rect 72660 3924 72666 3936
rect 74854 3924 74860 3936
rect 72660 3896 74860 3924
rect 72660 3884 72666 3896
rect 74854 3884 74860 3896
rect 74912 3884 74918 3936
rect 247630 3884 247636 3936
rect 247688 3924 247694 3936
rect 248598 3924 248604 3936
rect 247688 3896 248604 3924
rect 247688 3884 247694 3896
rect 248598 3884 248604 3896
rect 248656 3884 248662 3936
rect 285902 3884 285908 3936
rect 285960 3924 285966 3936
rect 287790 3924 287796 3936
rect 285960 3896 287796 3924
rect 285960 3884 285966 3896
rect 287790 3884 287796 3896
rect 287848 3884 287854 3936
rect 1670 3816 1676 3868
rect 1728 3856 1734 3868
rect 5210 3856 5216 3868
rect 1728 3828 5216 3856
rect 1728 3816 1734 3828
rect 5210 3816 5216 3828
rect 5268 3816 5274 3868
rect 13538 3816 13544 3868
rect 13596 3856 13602 3868
rect 16802 3856 16808 3868
rect 13596 3828 16808 3856
rect 13596 3816 13602 3828
rect 16802 3816 16808 3828
rect 16860 3816 16866 3868
rect 19426 3816 19432 3868
rect 19484 3856 19490 3868
rect 22598 3856 22604 3868
rect 19484 3828 22604 3856
rect 19484 3816 19490 3828
rect 22598 3816 22604 3828
rect 22656 3816 22662 3868
rect 23014 3816 23020 3868
rect 23072 3856 23078 3868
rect 26094 3856 26100 3868
rect 23072 3828 26100 3856
rect 23072 3816 23078 3828
rect 26094 3816 26100 3828
rect 26152 3816 26158 3868
rect 26510 3816 26516 3868
rect 26568 3856 26574 3868
rect 29590 3856 29596 3868
rect 26568 3828 29596 3856
rect 26568 3816 26574 3828
rect 29590 3816 29596 3828
rect 29648 3816 29654 3868
rect 30098 3816 30104 3868
rect 30156 3856 30162 3868
rect 33086 3856 33092 3868
rect 30156 3828 33092 3856
rect 30156 3816 30162 3828
rect 33086 3816 33092 3828
rect 33144 3816 33150 3868
rect 33594 3816 33600 3868
rect 33652 3856 33658 3868
rect 36582 3856 36588 3868
rect 33652 3828 36588 3856
rect 33652 3816 33658 3828
rect 36582 3816 36588 3828
rect 36640 3816 36646 3868
rect 37182 3816 37188 3868
rect 37240 3856 37246 3868
rect 39986 3856 39992 3868
rect 37240 3828 39992 3856
rect 37240 3816 37246 3828
rect 39986 3816 39992 3828
rect 40044 3816 40050 3868
rect 41874 3816 41880 3868
rect 41932 3856 41938 3868
rect 44678 3856 44684 3868
rect 41932 3828 44684 3856
rect 41932 3816 41938 3828
rect 44678 3816 44684 3828
rect 44736 3816 44742 3868
rect 45462 3816 45468 3868
rect 45520 3856 45526 3868
rect 48174 3856 48180 3868
rect 45520 3828 48180 3856
rect 45520 3816 45526 3828
rect 48174 3816 48180 3828
rect 48232 3816 48238 3868
rect 48958 3816 48964 3868
rect 49016 3856 49022 3868
rect 51578 3856 51584 3868
rect 49016 3828 51584 3856
rect 49016 3816 49022 3828
rect 51578 3816 51584 3828
rect 51636 3816 51642 3868
rect 53742 3816 53748 3868
rect 53800 3856 53806 3868
rect 56270 3856 56276 3868
rect 53800 3828 56276 3856
rect 53800 3816 53806 3828
rect 56270 3816 56276 3828
rect 56328 3816 56334 3868
rect 57238 3816 57244 3868
rect 57296 3856 57302 3868
rect 59766 3856 59772 3868
rect 57296 3828 59772 3856
rect 57296 3816 57302 3828
rect 59766 3816 59772 3828
rect 59824 3816 59830 3868
rect 71498 3816 71504 3868
rect 71556 3856 71562 3868
rect 73658 3856 73664 3868
rect 71556 3828 73664 3856
rect 71556 3816 71562 3828
rect 73658 3816 73664 3828
rect 73716 3816 73722 3868
rect 78582 3816 78588 3868
rect 78640 3856 78646 3868
rect 80650 3856 80656 3868
rect 78640 3828 80656 3856
rect 78640 3816 78646 3828
rect 80650 3816 80656 3828
rect 80708 3816 80714 3868
rect 80882 3816 80888 3868
rect 80940 3856 80946 3868
rect 82950 3856 82956 3868
rect 80940 3828 82956 3856
rect 80940 3816 80946 3828
rect 82950 3816 82956 3828
rect 83008 3816 83014 3868
rect 87966 3816 87972 3868
rect 88024 3856 88030 3868
rect 89942 3856 89948 3868
rect 88024 3828 89948 3856
rect 88024 3816 88030 3828
rect 89942 3816 89948 3828
rect 90000 3816 90006 3868
rect 96246 3816 96252 3868
rect 96304 3856 96310 3868
rect 98038 3856 98044 3868
rect 96304 3828 98044 3856
rect 96304 3816 96310 3828
rect 98038 3816 98044 3828
rect 98096 3816 98102 3868
rect 244134 3816 244140 3868
rect 244192 3856 244198 3868
rect 245194 3856 245200 3868
rect 244192 3828 245200 3856
rect 244192 3816 244198 3828
rect 245194 3816 245200 3828
rect 245252 3816 245258 3868
rect 256922 3816 256928 3868
rect 256980 3856 256986 3868
rect 258258 3856 258264 3868
rect 256980 3828 258264 3856
rect 256980 3816 256986 3828
rect 258258 3816 258264 3828
rect 258316 3816 258322 3868
rect 259222 3816 259228 3868
rect 259280 3856 259286 3868
rect 260650 3856 260656 3868
rect 259280 3828 260656 3856
rect 259280 3816 259286 3828
rect 260650 3816 260656 3828
rect 260708 3816 260714 3868
rect 261614 3816 261620 3868
rect 261672 3856 261678 3868
rect 262950 3856 262956 3868
rect 261672 3828 262956 3856
rect 261672 3816 261678 3828
rect 262950 3816 262956 3828
rect 263008 3816 263014 3868
rect 263914 3816 263920 3868
rect 263972 3856 263978 3868
rect 265342 3856 265348 3868
rect 263972 3828 265348 3856
rect 263972 3816 263978 3828
rect 265342 3816 265348 3828
rect 265400 3816 265406 3868
rect 268514 3816 268520 3868
rect 268572 3856 268578 3868
rect 270034 3856 270040 3868
rect 268572 3828 270040 3856
rect 268572 3816 268578 3828
rect 270034 3816 270040 3828
rect 270092 3816 270098 3868
rect 270814 3816 270820 3868
rect 270872 3856 270878 3868
rect 272426 3856 272432 3868
rect 270872 3828 272432 3856
rect 270872 3816 270878 3828
rect 272426 3816 272432 3828
rect 272484 3816 272490 3868
rect 275506 3816 275512 3868
rect 275564 3856 275570 3868
rect 277118 3856 277124 3868
rect 275564 3828 277124 3856
rect 275564 3816 275570 3828
rect 277118 3816 277124 3828
rect 277176 3816 277182 3868
rect 277806 3816 277812 3868
rect 277864 3856 277870 3868
rect 279510 3856 279516 3868
rect 277864 3828 279516 3856
rect 277864 3816 277870 3828
rect 279510 3816 279516 3828
rect 279568 3816 279574 3868
rect 284798 3816 284804 3868
rect 284856 3856 284862 3868
rect 286594 3856 286600 3868
rect 284856 3828 286600 3856
rect 284856 3816 284862 3828
rect 286594 3816 286600 3828
rect 286652 3816 286658 3868
rect 292894 3816 292900 3868
rect 292952 3856 292958 3868
rect 294874 3856 294880 3868
rect 292952 3828 294880 3856
rect 292952 3816 292958 3828
rect 294874 3816 294880 3828
rect 294932 3816 294938 3868
rect 299886 3816 299892 3868
rect 299944 3856 299950 3868
rect 301958 3856 301964 3868
rect 299944 3828 301964 3856
rect 299944 3816 299950 3828
rect 301958 3816 301964 3828
rect 302016 3816 302022 3868
rect 306786 3816 306792 3868
rect 306844 3856 306850 3868
rect 309042 3856 309048 3868
rect 306844 3828 309048 3856
rect 306844 3816 306850 3828
rect 309042 3816 309048 3828
rect 309100 3816 309106 3868
rect 566 3748 572 3800
rect 624 3788 630 3800
rect 4106 3788 4112 3800
rect 624 3760 4112 3788
rect 624 3748 630 3760
rect 4106 3748 4112 3760
rect 4164 3748 4170 3800
rect 7650 3748 7656 3800
rect 7708 3788 7714 3800
rect 11006 3788 11012 3800
rect 7708 3760 11012 3788
rect 7708 3748 7714 3760
rect 11006 3748 11012 3760
rect 11064 3748 11070 3800
rect 12342 3748 12348 3800
rect 12400 3788 12406 3800
rect 15698 3788 15704 3800
rect 12400 3760 15704 3788
rect 12400 3748 12406 3760
rect 15698 3748 15704 3760
rect 15756 3748 15762 3800
rect 15930 3748 15936 3800
rect 15988 3788 15994 3800
rect 19102 3788 19108 3800
rect 15988 3760 19108 3788
rect 15988 3748 15994 3760
rect 19102 3748 19108 3760
rect 19160 3748 19166 3800
rect 21818 3748 21824 3800
rect 21876 3788 21882 3800
rect 24898 3788 24904 3800
rect 21876 3760 24904 3788
rect 21876 3748 21882 3760
rect 24898 3748 24904 3760
rect 24956 3748 24962 3800
rect 25314 3748 25320 3800
rect 25372 3788 25378 3800
rect 28394 3788 28400 3800
rect 25372 3760 28400 3788
rect 25372 3748 25378 3760
rect 28394 3748 28400 3760
rect 28452 3748 28458 3800
rect 31294 3748 31300 3800
rect 31352 3788 31358 3800
rect 34190 3788 34196 3800
rect 31352 3760 34196 3788
rect 31352 3748 31358 3760
rect 34190 3748 34196 3760
rect 34248 3748 34254 3800
rect 34790 3748 34796 3800
rect 34848 3788 34854 3800
rect 37686 3788 37692 3800
rect 34848 3760 37692 3788
rect 34848 3748 34854 3760
rect 37686 3748 37692 3760
rect 37744 3748 37750 3800
rect 40678 3748 40684 3800
rect 40736 3788 40742 3800
rect 43482 3788 43488 3800
rect 40736 3760 43488 3788
rect 40736 3748 40742 3760
rect 43482 3748 43488 3760
rect 43540 3748 43546 3800
rect 44266 3748 44272 3800
rect 44324 3788 44330 3800
rect 46978 3788 46984 3800
rect 44324 3760 46984 3788
rect 44324 3748 44330 3760
rect 46978 3748 46984 3760
rect 47036 3748 47042 3800
rect 47854 3748 47860 3800
rect 47912 3788 47918 3800
rect 50474 3788 50480 3800
rect 47912 3760 50480 3788
rect 47912 3748 47918 3760
rect 50474 3748 50480 3760
rect 50532 3748 50538 3800
rect 51350 3748 51356 3800
rect 51408 3788 51414 3800
rect 53970 3788 53976 3800
rect 51408 3760 53976 3788
rect 51408 3748 51414 3760
rect 53970 3748 53976 3760
rect 54028 3748 54034 3800
rect 54938 3748 54944 3800
rect 54996 3788 55002 3800
rect 57374 3788 57380 3800
rect 54996 3760 57380 3788
rect 54996 3748 55002 3760
rect 57374 3748 57380 3760
rect 57432 3748 57438 3800
rect 58434 3748 58440 3800
rect 58492 3788 58498 3800
rect 60870 3788 60876 3800
rect 58492 3760 60876 3788
rect 58492 3748 58498 3760
rect 60870 3748 60876 3760
rect 60928 3748 60934 3800
rect 64322 3748 64328 3800
rect 64380 3788 64386 3800
rect 66666 3788 66672 3800
rect 64380 3760 66672 3788
rect 64380 3748 64386 3760
rect 66666 3748 66672 3760
rect 66724 3748 66730 3800
rect 67082 3748 67088 3800
rect 67140 3788 67146 3800
rect 69058 3788 69064 3800
rect 67140 3760 69064 3788
rect 67140 3748 67146 3760
rect 69058 3748 69064 3760
rect 69116 3748 69122 3800
rect 70302 3748 70308 3800
rect 70360 3788 70366 3800
rect 72462 3788 72468 3800
rect 70360 3760 72468 3788
rect 70360 3748 70366 3760
rect 72462 3748 72468 3760
rect 72520 3748 72526 3800
rect 73798 3748 73804 3800
rect 73856 3788 73862 3800
rect 75958 3788 75964 3800
rect 73856 3760 75964 3788
rect 73856 3748 73862 3760
rect 75958 3748 75964 3760
rect 76016 3748 76022 3800
rect 79686 3748 79692 3800
rect 79744 3788 79750 3800
rect 81754 3788 81760 3800
rect 79744 3760 81760 3788
rect 79744 3748 79750 3760
rect 81754 3748 81760 3760
rect 81812 3748 81818 3800
rect 86862 3748 86868 3800
rect 86920 3788 86926 3800
rect 88746 3788 88752 3800
rect 86920 3760 88752 3788
rect 86920 3748 86926 3760
rect 88746 3748 88752 3760
rect 88804 3748 88810 3800
rect 95142 3748 95148 3800
rect 95200 3788 95206 3800
rect 96842 3788 96848 3800
rect 95200 3760 96848 3788
rect 95200 3748 95206 3760
rect 96842 3748 96848 3760
rect 96900 3748 96906 3800
rect 103330 3748 103336 3800
rect 103388 3788 103394 3800
rect 104938 3788 104944 3800
rect 103388 3760 104944 3788
rect 103388 3748 103394 3760
rect 104938 3748 104944 3760
rect 104996 3748 105002 3800
rect 216350 3748 216356 3800
rect 216408 3788 216414 3800
rect 216858 3788 216864 3800
rect 216408 3760 216864 3788
rect 216408 3748 216414 3760
rect 216858 3748 216864 3760
rect 216916 3748 216922 3800
rect 222146 3748 222152 3800
rect 222204 3788 222210 3800
rect 222746 3788 222752 3800
rect 222204 3760 222752 3788
rect 222204 3748 222210 3760
rect 222746 3748 222752 3760
rect 222804 3748 222810 3800
rect 224446 3748 224452 3800
rect 224504 3788 224510 3800
rect 225138 3788 225144 3800
rect 224504 3760 225144 3788
rect 224504 3748 224510 3760
rect 225138 3748 225144 3760
rect 225196 3748 225202 3800
rect 230242 3748 230248 3800
rect 230300 3788 230306 3800
rect 231026 3788 231032 3800
rect 230300 3760 231032 3788
rect 230300 3748 230306 3760
rect 231026 3748 231032 3760
rect 231084 3748 231090 3800
rect 231438 3748 231444 3800
rect 231496 3788 231502 3800
rect 232222 3788 232228 3800
rect 231496 3760 232228 3788
rect 231496 3748 231502 3760
rect 232222 3748 232228 3760
rect 232280 3748 232286 3800
rect 232542 3748 232548 3800
rect 232600 3788 232606 3800
rect 233418 3788 233424 3800
rect 232600 3760 233424 3788
rect 232600 3748 232606 3760
rect 233418 3748 233424 3760
rect 233476 3748 233482 3800
rect 233738 3748 233744 3800
rect 233796 3788 233802 3800
rect 234614 3788 234620 3800
rect 233796 3760 234620 3788
rect 233796 3748 233802 3760
rect 234614 3748 234620 3760
rect 234672 3748 234678 3800
rect 237234 3748 237240 3800
rect 237292 3788 237298 3800
rect 238110 3788 238116 3800
rect 237292 3760 238116 3788
rect 237292 3748 237298 3760
rect 238110 3748 238116 3760
rect 238168 3748 238174 3800
rect 238338 3748 238344 3800
rect 238396 3788 238402 3800
rect 239306 3788 239312 3800
rect 238396 3760 239312 3788
rect 238396 3748 238402 3760
rect 239306 3748 239312 3760
rect 239364 3748 239370 3800
rect 239534 3748 239540 3800
rect 239592 3788 239598 3800
rect 240502 3788 240508 3800
rect 239592 3760 240508 3788
rect 239592 3748 239598 3760
rect 240502 3748 240508 3760
rect 240560 3748 240566 3800
rect 240730 3748 240736 3800
rect 240788 3788 240794 3800
rect 241698 3788 241704 3800
rect 240788 3760 241704 3788
rect 240788 3748 240794 3760
rect 241698 3748 241704 3760
rect 241756 3748 241762 3800
rect 241834 3748 241840 3800
rect 241892 3788 241898 3800
rect 242894 3788 242900 3800
rect 241892 3760 242900 3788
rect 241892 3748 241898 3760
rect 242894 3748 242900 3760
rect 242952 3748 242958 3800
rect 245330 3748 245336 3800
rect 245388 3788 245394 3800
rect 246390 3788 246396 3800
rect 245388 3760 246396 3788
rect 245388 3748 245394 3760
rect 246390 3748 246396 3760
rect 246448 3748 246454 3800
rect 246526 3748 246532 3800
rect 246584 3788 246590 3800
rect 247586 3788 247592 3800
rect 246584 3760 247592 3788
rect 246584 3748 246590 3760
rect 247586 3748 247592 3760
rect 247644 3748 247650 3800
rect 250022 3748 250028 3800
rect 250080 3788 250086 3800
rect 251174 3788 251180 3800
rect 250080 3760 251180 3788
rect 250080 3748 250086 3760
rect 251174 3748 251180 3760
rect 251232 3748 251238 3800
rect 252322 3748 252328 3800
rect 252380 3788 252386 3800
rect 253474 3788 253480 3800
rect 252380 3760 253480 3788
rect 252380 3748 252386 3760
rect 253474 3748 253480 3760
rect 253532 3748 253538 3800
rect 255818 3748 255824 3800
rect 255876 3788 255882 3800
rect 257062 3788 257068 3800
rect 255876 3760 257068 3788
rect 255876 3748 255882 3760
rect 257062 3748 257068 3760
rect 257120 3748 257126 3800
rect 258118 3748 258124 3800
rect 258176 3788 258182 3800
rect 259454 3788 259460 3800
rect 258176 3760 259460 3788
rect 258176 3748 258182 3760
rect 259454 3748 259460 3760
rect 259512 3748 259518 3800
rect 260418 3748 260424 3800
rect 260476 3788 260482 3800
rect 261754 3788 261760 3800
rect 260476 3760 261760 3788
rect 260476 3748 260482 3760
rect 261754 3748 261760 3760
rect 261812 3748 261818 3800
rect 262718 3748 262724 3800
rect 262776 3788 262782 3800
rect 264146 3788 264152 3800
rect 262776 3760 264152 3788
rect 262776 3748 262782 3760
rect 264146 3748 264152 3760
rect 264204 3748 264210 3800
rect 265018 3748 265024 3800
rect 265076 3788 265082 3800
rect 266538 3788 266544 3800
rect 265076 3760 266544 3788
rect 265076 3748 265082 3760
rect 266538 3748 266544 3760
rect 266596 3748 266602 3800
rect 267410 3748 267416 3800
rect 267468 3788 267474 3800
rect 268838 3788 268844 3800
rect 267468 3760 268844 3788
rect 267468 3748 267474 3760
rect 268838 3748 268844 3760
rect 268896 3748 268902 3800
rect 269710 3748 269716 3800
rect 269768 3788 269774 3800
rect 271230 3788 271236 3800
rect 269768 3760 271236 3788
rect 269768 3748 269774 3760
rect 271230 3748 271236 3760
rect 271288 3748 271294 3800
rect 272010 3748 272016 3800
rect 272068 3788 272074 3800
rect 273622 3788 273628 3800
rect 272068 3760 273628 3788
rect 272068 3748 272074 3760
rect 273622 3748 273628 3760
rect 273680 3748 273686 3800
rect 276702 3748 276708 3800
rect 276760 3788 276766 3800
rect 278314 3788 278320 3800
rect 276760 3760 278320 3788
rect 276760 3748 276766 3760
rect 278314 3748 278320 3760
rect 278372 3748 278378 3800
rect 279002 3748 279008 3800
rect 279060 3788 279066 3800
rect 280706 3788 280712 3800
rect 279060 3760 280712 3788
rect 279060 3748 279066 3760
rect 280706 3748 280712 3760
rect 280764 3748 280770 3800
rect 283602 3748 283608 3800
rect 283660 3788 283666 3800
rect 285398 3788 285404 3800
rect 283660 3760 285404 3788
rect 283660 3748 283666 3760
rect 285398 3748 285404 3760
rect 285456 3748 285462 3800
rect 287098 3748 287104 3800
rect 287156 3788 287162 3800
rect 288986 3788 288992 3800
rect 287156 3760 288992 3788
rect 287156 3748 287162 3760
rect 288986 3748 288992 3760
rect 289044 3748 289050 3800
rect 291698 3748 291704 3800
rect 291756 3788 291762 3800
rect 293678 3788 293684 3800
rect 291756 3760 293684 3788
rect 291756 3748 291762 3760
rect 293678 3748 293684 3760
rect 293736 3748 293742 3800
rect 294090 3748 294096 3800
rect 294148 3788 294154 3800
rect 296070 3788 296076 3800
rect 294148 3760 296076 3788
rect 294148 3748 294154 3760
rect 296070 3748 296076 3760
rect 296128 3748 296134 3800
rect 298690 3748 298696 3800
rect 298748 3788 298754 3800
rect 300762 3788 300768 3800
rect 298748 3760 300768 3788
rect 298748 3748 298754 3760
rect 300762 3748 300768 3760
rect 300820 3748 300826 3800
rect 300990 3748 300996 3800
rect 301048 3788 301054 3800
rect 303154 3788 303160 3800
rect 301048 3760 303160 3788
rect 301048 3748 301054 3760
rect 303154 3748 303160 3760
rect 303212 3748 303218 3800
rect 307982 3748 307988 3800
rect 308040 3788 308046 3800
rect 310238 3788 310244 3800
rect 308040 3760 310244 3788
rect 308040 3748 308046 3760
rect 310238 3748 310244 3760
rect 310296 3748 310302 3800
rect 316078 3748 316084 3800
rect 316136 3788 316142 3800
rect 318518 3788 318524 3800
rect 316136 3760 318524 3788
rect 316136 3748 316142 3760
rect 318518 3748 318524 3760
rect 318576 3748 318582 3800
rect 323070 3748 323076 3800
rect 323128 3788 323134 3800
rect 325602 3788 325608 3800
rect 323128 3760 325608 3788
rect 323128 3748 323134 3760
rect 325602 3748 325608 3760
rect 325660 3748 325666 3800
rect 6454 3000 6460 3052
rect 6512 3040 6518 3052
rect 9858 3040 9864 3052
rect 6512 3012 9864 3040
rect 6512 3000 6518 3012
rect 9858 3000 9864 3012
rect 9916 3000 9922 3052
rect 63218 3000 63224 3052
rect 63276 3040 63282 3052
rect 65518 3040 65524 3052
rect 63276 3012 65524 3040
rect 63276 3000 63282 3012
rect 65518 3000 65524 3012
rect 65576 3000 65582 3052
rect 535362 2932 535368 2984
rect 535420 2972 535426 2984
rect 541986 2972 541992 2984
rect 535420 2944 541992 2972
rect 535420 2932 535426 2944
rect 541986 2932 541992 2944
rect 542044 2932 542050 2984
rect 573634 2932 573640 2984
rect 573692 2972 573698 2984
rect 580994 2972 581000 2984
rect 573692 2944 581000 2972
rect 573692 2932 573698 2944
rect 580994 2932 581000 2944
rect 581052 2932 581058 2984
rect 18230 2864 18236 2916
rect 18288 2904 18294 2916
rect 21450 2904 21456 2916
rect 18288 2876 21456 2904
rect 18288 2864 18294 2876
rect 21450 2864 21456 2876
rect 21508 2864 21514 2916
rect 253382 2864 253388 2916
rect 253440 2904 253446 2916
rect 254670 2904 254676 2916
rect 253440 2876 254676 2904
rect 253440 2864 253446 2876
rect 254670 2864 254676 2876
rect 254728 2864 254734 2916
rect 506382 2864 506388 2916
rect 506440 2904 506446 2916
rect 512454 2904 512460 2916
rect 506440 2876 512460 2904
rect 506440 2864 506446 2876
rect 512454 2864 512460 2876
rect 512512 2864 512518 2916
rect 516778 2864 516784 2916
rect 516836 2904 516842 2916
rect 523034 2904 523040 2916
rect 516836 2876 523040 2904
rect 516836 2864 516842 2876
rect 523034 2864 523040 2876
rect 523092 2864 523098 2916
rect 524966 2864 524972 2916
rect 525024 2904 525030 2916
rect 531314 2904 531320 2916
rect 525024 2876 531320 2904
rect 525024 2864 525030 2876
rect 531314 2864 531320 2876
rect 531372 2864 531378 2916
rect 536558 2864 536564 2916
rect 536616 2904 536622 2916
rect 543182 2904 543188 2916
rect 536616 2876 543188 2904
rect 536616 2864 536622 2876
rect 543182 2864 543188 2876
rect 543240 2864 543246 2916
rect 544654 2864 544660 2916
rect 544712 2904 544718 2916
rect 551462 2904 551468 2916
rect 544712 2876 551468 2904
rect 544712 2864 544718 2876
rect 551462 2864 551468 2876
rect 551520 2864 551526 2916
rect 553946 2864 553952 2916
rect 554004 2904 554010 2916
rect 560846 2904 560852 2916
rect 554004 2876 560852 2904
rect 554004 2864 554010 2876
rect 560846 2864 560852 2876
rect 560904 2864 560910 2916
rect 574830 2864 574836 2916
rect 574888 2904 574894 2916
rect 582190 2904 582196 2916
rect 574888 2876 582196 2904
rect 574888 2864 574894 2876
rect 582190 2864 582196 2876
rect 582248 2864 582254 2916
rect 4062 2796 4068 2848
rect 4120 2836 4126 2848
rect 7466 2836 7472 2848
rect 4120 2808 7472 2836
rect 4120 2796 4126 2808
rect 7466 2796 7472 2808
rect 7524 2796 7530 2848
rect 9950 2796 9956 2848
rect 10008 2836 10014 2848
rect 13262 2836 13268 2848
rect 10008 2808 13268 2836
rect 10008 2796 10014 2808
rect 13262 2796 13268 2808
rect 13320 2796 13326 2848
rect 17034 2796 17040 2848
rect 17092 2836 17098 2848
rect 20254 2836 20260 2848
rect 17092 2808 20260 2836
rect 17092 2796 17098 2808
rect 20254 2796 20260 2808
rect 20312 2796 20318 2848
rect 28902 2796 28908 2848
rect 28960 2836 28966 2848
rect 31846 2836 31852 2848
rect 28960 2808 31852 2836
rect 28960 2796 28966 2808
rect 31846 2796 31852 2808
rect 31904 2796 31910 2848
rect 35986 2796 35992 2848
rect 36044 2836 36050 2848
rect 38838 2836 38844 2848
rect 36044 2808 38844 2836
rect 36044 2796 36050 2808
rect 38838 2796 38844 2808
rect 38896 2796 38902 2848
rect 39574 2796 39580 2848
rect 39632 2836 39638 2848
rect 42334 2836 42340 2848
rect 39632 2808 42340 2836
rect 39632 2796 39638 2808
rect 42334 2796 42340 2808
rect 42392 2796 42398 2848
rect 62022 2796 62028 2848
rect 62080 2836 62086 2848
rect 64414 2836 64420 2848
rect 62080 2808 64420 2836
rect 62080 2796 62086 2808
rect 64414 2796 64420 2808
rect 64472 2796 64478 2848
rect 65518 2796 65524 2848
rect 65576 2836 65582 2848
rect 67818 2836 67824 2848
rect 65576 2808 67824 2836
rect 65576 2796 65582 2808
rect 67818 2796 67824 2808
rect 67876 2796 67882 2848
rect 248874 2796 248880 2848
rect 248932 2836 248938 2848
rect 249978 2836 249984 2848
rect 248932 2808 249984 2836
rect 248932 2796 248938 2808
rect 249978 2796 249984 2808
rect 250036 2796 250042 2848
rect 251082 2796 251088 2848
rect 251140 2836 251146 2848
rect 252370 2836 252376 2848
rect 251140 2808 252376 2836
rect 251140 2796 251146 2808
rect 252370 2796 252376 2808
rect 252428 2796 252434 2848
rect 254578 2796 254584 2848
rect 254636 2836 254642 2848
rect 255866 2836 255872 2848
rect 254636 2808 255872 2836
rect 254636 2796 254642 2808
rect 255866 2796 255872 2808
rect 255924 2796 255930 2848
rect 309226 2796 309232 2848
rect 309284 2836 309290 2848
rect 311434 2836 311440 2848
rect 309284 2808 311440 2836
rect 309284 2796 309290 2808
rect 311434 2796 311440 2808
rect 311492 2796 311498 2848
rect 315022 2796 315028 2848
rect 315080 2836 315086 2848
rect 317322 2836 317328 2848
rect 315080 2808 317328 2836
rect 315080 2796 315086 2808
rect 317322 2796 317328 2808
rect 317380 2796 317386 2848
rect 411162 2796 411168 2848
rect 411220 2836 411226 2848
rect 415486 2836 415492 2848
rect 411220 2808 415492 2836
rect 411220 2796 411226 2808
rect 415486 2796 415492 2808
rect 415544 2796 415550 2848
rect 440142 2796 440148 2848
rect 440200 2836 440206 2848
rect 445018 2836 445024 2848
rect 440200 2808 445024 2836
rect 440200 2796 440206 2808
rect 445018 2796 445024 2808
rect 445076 2796 445082 2848
rect 449526 2796 449532 2848
rect 449584 2836 449590 2848
rect 454494 2836 454500 2848
rect 449584 2808 454500 2836
rect 449584 2796 449590 2808
rect 454494 2796 454500 2808
rect 454552 2796 454558 2848
rect 478506 2796 478512 2848
rect 478564 2836 478570 2848
rect 484026 2836 484032 2848
rect 478564 2808 484032 2836
rect 478564 2796 478570 2808
rect 484026 2796 484032 2808
rect 484084 2796 484090 2848
rect 487798 2796 487804 2848
rect 487856 2836 487862 2848
rect 493502 2836 493508 2848
rect 487856 2808 493508 2836
rect 487856 2796 487862 2808
rect 493502 2796 493508 2808
rect 493560 2796 493566 2848
rect 507578 2796 507584 2848
rect 507636 2836 507642 2848
rect 513558 2836 513564 2848
rect 507636 2808 513564 2836
rect 507636 2796 507642 2808
rect 513558 2796 513564 2808
rect 513616 2796 513622 2848
rect 515674 2796 515680 2848
rect 515732 2836 515738 2848
rect 521838 2836 521844 2848
rect 515732 2808 521844 2836
rect 515732 2796 515738 2808
rect 521838 2796 521844 2808
rect 521896 2796 521902 2848
rect 545850 2796 545856 2848
rect 545908 2836 545914 2848
rect 552658 2836 552664 2848
rect 545908 2808 552664 2836
rect 545908 2796 545914 2808
rect 552658 2796 552664 2808
rect 552716 2796 552722 2848
rect 3234 1300 3240 1352
rect 3292 1340 3298 1352
rect 6362 1340 6368 1352
rect 3292 1312 6368 1340
rect 3292 1300 3298 1312
rect 6362 1300 6368 1312
rect 6420 1300 6426 1352
rect 60826 1300 60832 1352
rect 60884 1340 60890 1352
rect 63310 1340 63316 1352
rect 60884 1312 63316 1340
rect 60884 1300 60890 1312
rect 63310 1300 63316 1312
rect 63368 1300 63374 1352
rect 67910 1300 67916 1352
rect 67968 1340 67974 1352
rect 70118 1340 70124 1352
rect 67968 1312 70124 1340
rect 67968 1300 67974 1312
rect 70118 1300 70124 1312
rect 70176 1300 70182 1352
rect 76190 1300 76196 1352
rect 76248 1340 76254 1352
rect 78214 1340 78220 1352
rect 76248 1312 78220 1340
rect 76248 1300 76254 1312
rect 78214 1300 78220 1312
rect 78272 1300 78278 1352
rect 83274 1300 83280 1352
rect 83332 1340 83338 1352
rect 85206 1340 85212 1352
rect 83332 1312 85212 1340
rect 83332 1300 83338 1312
rect 85206 1300 85212 1312
rect 85264 1300 85270 1352
rect 85666 1300 85672 1352
rect 85724 1340 85730 1352
rect 87506 1340 87512 1352
rect 85724 1312 87512 1340
rect 85724 1300 85730 1312
rect 87506 1300 87512 1312
rect 87564 1300 87570 1352
rect 89162 1300 89168 1352
rect 89220 1340 89226 1352
rect 91002 1340 91008 1352
rect 89220 1312 91008 1340
rect 89220 1300 89226 1312
rect 91002 1300 91008 1312
rect 91060 1300 91066 1352
rect 91554 1300 91560 1352
rect 91612 1340 91618 1352
rect 93302 1340 93308 1352
rect 91612 1312 93308 1340
rect 91612 1300 91618 1312
rect 93302 1300 93308 1312
rect 93360 1300 93366 1352
rect 93946 1300 93952 1352
rect 94004 1340 94010 1352
rect 95694 1340 95700 1352
rect 94004 1312 95700 1340
rect 94004 1300 94010 1312
rect 95694 1300 95700 1312
rect 95752 1300 95758 1352
rect 97442 1300 97448 1352
rect 97500 1340 97506 1352
rect 99098 1340 99104 1352
rect 97500 1312 99104 1340
rect 97500 1300 97506 1312
rect 99098 1300 99104 1312
rect 99156 1300 99162 1352
rect 101030 1300 101036 1352
rect 101088 1340 101094 1352
rect 102594 1340 102600 1352
rect 101088 1312 102600 1340
rect 101088 1300 101094 1312
rect 102594 1300 102600 1312
rect 102652 1300 102658 1352
rect 104526 1300 104532 1352
rect 104584 1340 104590 1352
rect 106090 1340 106096 1352
rect 104584 1312 106096 1340
rect 104584 1300 104590 1312
rect 106090 1300 106096 1312
rect 106148 1300 106154 1352
rect 106918 1300 106924 1352
rect 106976 1340 106982 1352
rect 108390 1340 108396 1352
rect 106976 1312 108396 1340
rect 106976 1300 106982 1312
rect 108390 1300 108396 1312
rect 108448 1300 108454 1352
rect 109310 1300 109316 1352
rect 109368 1340 109374 1352
rect 110690 1340 110696 1352
rect 109368 1312 110696 1340
rect 109368 1300 109374 1312
rect 110690 1300 110696 1312
rect 110748 1300 110754 1352
rect 112806 1300 112812 1352
rect 112864 1340 112870 1352
rect 114186 1340 114192 1352
rect 112864 1312 114192 1340
rect 112864 1300 112870 1312
rect 114186 1300 114192 1312
rect 114244 1300 114250 1352
rect 116394 1300 116400 1352
rect 116452 1340 116458 1352
rect 117682 1340 117688 1352
rect 116452 1312 117688 1340
rect 116452 1300 116458 1312
rect 117682 1300 117688 1312
rect 117740 1300 117746 1352
rect 119890 1300 119896 1352
rect 119948 1340 119954 1352
rect 121178 1340 121184 1352
rect 119948 1312 121184 1340
rect 119948 1300 119954 1312
rect 121178 1300 121184 1312
rect 121236 1300 121242 1352
rect 125870 1300 125876 1352
rect 125928 1340 125934 1352
rect 126974 1340 126980 1352
rect 125928 1312 126980 1340
rect 125928 1300 125934 1312
rect 126974 1300 126980 1312
rect 127032 1300 127038 1352
rect 129366 1300 129372 1352
rect 129424 1340 129430 1352
rect 130470 1340 130476 1352
rect 129424 1312 130476 1340
rect 129424 1300 129430 1312
rect 130470 1300 130476 1312
rect 130528 1300 130534 1352
rect 130562 1300 130568 1352
rect 130620 1340 130626 1352
rect 131574 1340 131580 1352
rect 130620 1312 131580 1340
rect 130620 1300 130626 1312
rect 131574 1300 131580 1312
rect 131632 1300 131638 1352
rect 131758 1300 131764 1352
rect 131816 1340 131822 1352
rect 132770 1340 132776 1352
rect 131816 1312 132776 1340
rect 131816 1300 131822 1312
rect 132770 1300 132776 1312
rect 132828 1300 132834 1352
rect 132954 1300 132960 1352
rect 133012 1340 133018 1352
rect 133966 1340 133972 1352
rect 133012 1312 133972 1340
rect 133012 1300 133018 1312
rect 133966 1300 133972 1312
rect 134024 1300 134030 1352
rect 137646 1300 137652 1352
rect 137704 1340 137710 1352
rect 138566 1340 138572 1352
rect 137704 1312 138572 1340
rect 137704 1300 137710 1312
rect 138566 1300 138572 1312
rect 138624 1300 138630 1352
rect 144730 1300 144736 1352
rect 144788 1340 144794 1352
rect 145558 1340 145564 1352
rect 144788 1312 145564 1340
rect 144788 1300 144794 1312
rect 145558 1300 145564 1312
rect 145616 1300 145622 1352
rect 145926 1300 145932 1352
rect 145984 1340 145990 1352
rect 146662 1340 146668 1352
rect 145984 1312 146668 1340
rect 145984 1300 145990 1312
rect 146662 1300 146668 1312
rect 146720 1300 146726 1352
rect 148318 1300 148324 1352
rect 148376 1340 148382 1352
rect 149054 1340 149060 1352
rect 148376 1312 149060 1340
rect 148376 1300 148382 1312
rect 149054 1300 149060 1312
rect 149112 1300 149118 1352
rect 154206 1300 154212 1352
rect 154264 1340 154270 1352
rect 154850 1340 154856 1352
rect 154264 1312 154856 1340
rect 154264 1300 154270 1312
rect 154850 1300 154856 1312
rect 154908 1300 154914 1352
rect 162486 1300 162492 1352
rect 162544 1340 162550 1352
rect 162946 1340 162952 1352
rect 162544 1312 162952 1340
rect 162544 1300 162550 1312
rect 162946 1300 162952 1312
rect 163004 1300 163010 1352
rect 266262 1300 266268 1352
rect 266320 1340 266326 1352
rect 267734 1340 267740 1352
rect 266320 1312 267740 1340
rect 266320 1300 266326 1312
rect 267734 1300 267740 1312
rect 267792 1300 267798 1352
rect 273162 1300 273168 1352
rect 273220 1340 273226 1352
rect 274818 1340 274824 1352
rect 273220 1312 274824 1340
rect 273220 1300 273226 1312
rect 274818 1300 274824 1312
rect 274876 1300 274882 1352
rect 280062 1300 280068 1352
rect 280120 1340 280126 1352
rect 281902 1340 281908 1352
rect 280120 1312 281908 1340
rect 280120 1300 280126 1312
rect 281902 1300 281908 1312
rect 281960 1300 281966 1352
rect 282546 1300 282552 1352
rect 282604 1340 282610 1352
rect 284294 1340 284300 1352
rect 282604 1312 284300 1340
rect 282604 1300 282610 1312
rect 284294 1300 284300 1312
rect 284352 1300 284358 1352
rect 288342 1300 288348 1352
rect 288400 1340 288406 1352
rect 290182 1340 290188 1352
rect 288400 1312 290188 1340
rect 288400 1300 288406 1312
rect 290182 1300 290188 1312
rect 290240 1300 290246 1352
rect 295242 1300 295248 1352
rect 295300 1340 295306 1352
rect 297266 1340 297272 1352
rect 295300 1312 297272 1340
rect 295300 1300 295306 1312
rect 297266 1300 297272 1312
rect 297324 1300 297330 1352
rect 297542 1300 297548 1352
rect 297600 1340 297606 1352
rect 299658 1340 299664 1352
rect 297600 1312 299664 1340
rect 297600 1300 297606 1312
rect 299658 1300 299664 1312
rect 299716 1300 299722 1352
rect 302142 1300 302148 1352
rect 302200 1340 302206 1352
rect 304350 1340 304356 1352
rect 302200 1312 304356 1340
rect 302200 1300 302206 1312
rect 304350 1300 304356 1312
rect 304408 1300 304414 1352
rect 305730 1300 305736 1352
rect 305788 1340 305794 1352
rect 307938 1340 307944 1352
rect 305788 1312 307944 1340
rect 305788 1300 305794 1312
rect 307938 1300 307944 1312
rect 307996 1300 308002 1352
rect 310330 1300 310336 1352
rect 310388 1340 310394 1352
rect 312630 1340 312636 1352
rect 310388 1312 312636 1340
rect 310388 1300 310394 1312
rect 312630 1300 312636 1312
rect 312688 1300 312694 1352
rect 313826 1300 313832 1352
rect 313884 1340 313890 1352
rect 316218 1340 316224 1352
rect 313884 1312 316224 1340
rect 313884 1300 313890 1312
rect 316218 1300 316224 1312
rect 316276 1300 316282 1352
rect 317230 1300 317236 1352
rect 317288 1340 317294 1352
rect 319714 1340 319720 1352
rect 317288 1312 319720 1340
rect 317288 1300 317294 1312
rect 319714 1300 319720 1312
rect 319772 1300 319778 1352
rect 321922 1300 321928 1352
rect 321980 1340 321986 1352
rect 324406 1340 324412 1352
rect 321980 1312 324412 1340
rect 321980 1300 321986 1312
rect 324406 1300 324412 1312
rect 324464 1300 324470 1352
rect 325418 1300 325424 1352
rect 325476 1340 325482 1352
rect 327994 1340 328000 1352
rect 325476 1312 328000 1340
rect 325476 1300 325482 1312
rect 327994 1300 328000 1312
rect 328052 1300 328058 1352
rect 328914 1300 328920 1352
rect 328972 1340 328978 1352
rect 331582 1340 331588 1352
rect 328972 1312 331588 1340
rect 328972 1300 328978 1312
rect 331582 1300 331588 1312
rect 331640 1300 331646 1352
rect 332410 1300 332416 1352
rect 332468 1340 332474 1352
rect 335078 1340 335084 1352
rect 332468 1312 335084 1340
rect 332468 1300 332474 1312
rect 335078 1300 335084 1312
rect 335136 1300 335142 1352
rect 335906 1300 335912 1352
rect 335964 1340 335970 1352
rect 338666 1340 338672 1352
rect 335964 1312 338672 1340
rect 335964 1300 335970 1312
rect 338666 1300 338672 1312
rect 338724 1300 338730 1352
rect 339310 1300 339316 1352
rect 339368 1340 339374 1352
rect 342162 1340 342168 1352
rect 339368 1312 342168 1340
rect 339368 1300 339374 1312
rect 342162 1300 342168 1312
rect 342220 1300 342226 1352
rect 345106 1300 345112 1352
rect 345164 1340 345170 1352
rect 348050 1340 348056 1352
rect 345164 1312 348056 1340
rect 345164 1300 345170 1312
rect 348050 1300 348056 1312
rect 348108 1300 348114 1352
rect 349798 1300 349804 1352
rect 349856 1340 349862 1352
rect 352834 1340 352840 1352
rect 349856 1312 352840 1340
rect 349856 1300 349862 1312
rect 352834 1300 352840 1312
rect 352892 1300 352898 1352
rect 353202 1300 353208 1352
rect 353260 1340 353266 1352
rect 356330 1340 356336 1352
rect 353260 1312 356336 1340
rect 353260 1300 353266 1312
rect 356330 1300 356336 1312
rect 356388 1300 356394 1352
rect 356698 1300 356704 1352
rect 356756 1340 356762 1352
rect 359918 1340 359924 1352
rect 356756 1312 359924 1340
rect 356756 1300 356762 1312
rect 359918 1300 359924 1312
rect 359976 1300 359982 1352
rect 362586 1300 362592 1352
rect 362644 1340 362650 1352
rect 365806 1340 365812 1352
rect 362644 1312 365812 1340
rect 362644 1300 362650 1312
rect 365806 1300 365812 1312
rect 365864 1300 365870 1352
rect 367186 1300 367192 1352
rect 367244 1340 367250 1352
rect 370590 1340 370596 1352
rect 367244 1312 370596 1340
rect 367244 1300 367250 1312
rect 370590 1300 370596 1312
rect 370648 1300 370654 1352
rect 370682 1300 370688 1352
rect 370740 1340 370746 1352
rect 374086 1340 374092 1352
rect 370740 1312 374092 1340
rect 370740 1300 370746 1312
rect 374086 1300 374092 1312
rect 374144 1300 374150 1352
rect 376386 1300 376392 1352
rect 376444 1340 376450 1352
rect 379974 1340 379980 1352
rect 376444 1312 379980 1340
rect 376444 1300 376450 1312
rect 379974 1300 379980 1312
rect 380032 1300 380038 1352
rect 385770 1300 385776 1352
rect 385828 1340 385834 1352
rect 389450 1340 389456 1352
rect 385828 1312 389456 1340
rect 385828 1300 385834 1312
rect 389450 1300 389456 1312
rect 389508 1300 389514 1352
rect 395062 1300 395068 1352
rect 395120 1340 395126 1352
rect 398926 1340 398932 1352
rect 395120 1312 398932 1340
rect 395120 1300 395126 1312
rect 398926 1300 398932 1312
rect 398984 1300 398990 1352
rect 399662 1300 399668 1352
rect 399720 1340 399726 1352
rect 403618 1340 403624 1352
rect 399720 1312 403624 1340
rect 399720 1300 399726 1312
rect 403618 1300 403624 1312
rect 403676 1300 403682 1352
rect 405458 1300 405464 1352
rect 405516 1340 405522 1352
rect 409598 1340 409604 1352
rect 405516 1312 409604 1340
rect 405516 1300 405522 1312
rect 409598 1300 409604 1312
rect 409656 1300 409662 1352
rect 413554 1300 413560 1352
rect 413612 1340 413618 1352
rect 417878 1340 417884 1352
rect 413612 1312 417884 1340
rect 413612 1300 413618 1312
rect 417878 1300 417884 1312
rect 417936 1300 417942 1352
rect 422846 1300 422852 1352
rect 422904 1340 422910 1352
rect 427262 1340 427268 1352
rect 422904 1312 427268 1340
rect 422904 1300 422910 1312
rect 427262 1300 427268 1312
rect 427320 1300 427326 1352
rect 427538 1300 427544 1352
rect 427596 1340 427602 1352
rect 431862 1340 431868 1352
rect 427596 1312 431868 1340
rect 427596 1300 427602 1312
rect 431862 1300 431868 1312
rect 431920 1300 431926 1352
rect 433242 1300 433248 1352
rect 433300 1340 433306 1352
rect 437842 1340 437848 1352
rect 433300 1312 437848 1340
rect 433300 1300 433306 1312
rect 437842 1300 437848 1312
rect 437900 1300 437906 1352
rect 442626 1300 442632 1352
rect 442684 1340 442690 1352
rect 447410 1340 447416 1352
rect 442684 1312 447416 1340
rect 442684 1300 442690 1312
rect 447410 1300 447416 1312
rect 447468 1300 447474 1352
rect 448422 1300 448428 1352
rect 448480 1340 448486 1352
rect 453298 1340 453304 1352
rect 448480 1312 453304 1340
rect 448480 1300 448486 1312
rect 453298 1300 453304 1312
rect 453356 1300 453362 1352
rect 458818 1300 458824 1352
rect 458876 1340 458882 1352
rect 463970 1340 463976 1352
rect 458876 1312 463976 1340
rect 458876 1300 458882 1312
rect 463970 1300 463976 1312
rect 464028 1300 464034 1352
rect 468110 1300 468116 1352
rect 468168 1340 468174 1352
rect 473078 1340 473084 1352
rect 468168 1312 473084 1340
rect 468168 1300 468174 1312
rect 473078 1300 473084 1312
rect 473136 1300 473142 1352
rect 475102 1300 475108 1352
rect 475160 1340 475166 1352
rect 480530 1340 480536 1352
rect 475160 1312 480536 1340
rect 475160 1300 475166 1312
rect 480530 1300 480536 1312
rect 480588 1300 480594 1352
rect 485498 1300 485504 1352
rect 485556 1340 485562 1352
rect 490742 1340 490748 1352
rect 485556 1312 490748 1340
rect 485556 1300 485562 1312
rect 490742 1300 490748 1312
rect 490800 1300 490806 1352
rect 497090 1300 497096 1352
rect 497148 1340 497154 1352
rect 502978 1340 502984 1352
rect 497148 1312 502984 1340
rect 497148 1300 497154 1312
rect 502978 1300 502984 1312
rect 503036 1300 503042 1352
rect 504082 1300 504088 1352
rect 504140 1340 504146 1352
rect 509694 1340 509700 1352
rect 504140 1312 509700 1340
rect 504140 1300 504146 1312
rect 509694 1300 509700 1312
rect 509752 1300 509758 1352
rect 513282 1300 513288 1352
rect 513340 1340 513346 1352
rect 519538 1340 519544 1352
rect 513340 1312 519544 1340
rect 513340 1300 513346 1312
rect 519538 1300 519544 1312
rect 519596 1300 519602 1352
rect 526070 1300 526076 1352
rect 526128 1340 526134 1352
rect 532142 1340 532148 1352
rect 526128 1312 532148 1340
rect 526128 1300 526134 1312
rect 532142 1300 532148 1312
rect 532200 1300 532206 1352
rect 534258 1300 534264 1352
rect 534316 1340 534322 1352
rect 540422 1340 540428 1352
rect 534316 1312 540428 1340
rect 534316 1300 534322 1312
rect 540422 1300 540428 1312
rect 540480 1300 540486 1352
rect 541158 1300 541164 1352
rect 541216 1340 541222 1352
rect 547874 1340 547880 1352
rect 541216 1312 547880 1340
rect 541216 1300 541222 1312
rect 547874 1300 547880 1312
rect 547932 1300 547938 1352
rect 548150 1300 548156 1352
rect 548208 1340 548214 1352
rect 554774 1340 554780 1352
rect 548208 1312 554780 1340
rect 548208 1300 548214 1312
rect 554774 1300 554780 1312
rect 554832 1300 554838 1352
rect 555142 1300 555148 1352
rect 555200 1340 555206 1352
rect 562042 1340 562048 1352
rect 555200 1312 562048 1340
rect 555200 1300 555206 1312
rect 562042 1300 562048 1312
rect 562100 1300 562106 1352
rect 566734 1300 566740 1352
rect 566792 1340 566798 1352
rect 566792 1312 571288 1340
rect 566792 1300 566798 1312
rect 74994 1232 75000 1284
rect 75052 1272 75058 1284
rect 77110 1272 77116 1284
rect 75052 1244 77116 1272
rect 75052 1232 75058 1244
rect 77110 1232 77116 1244
rect 77168 1232 77174 1284
rect 77386 1232 77392 1284
rect 77444 1272 77450 1284
rect 79410 1272 79416 1284
rect 77444 1244 79416 1272
rect 77444 1232 77450 1244
rect 79410 1232 79416 1244
rect 79468 1232 79474 1284
rect 82078 1232 82084 1284
rect 82136 1272 82142 1284
rect 84010 1272 84016 1284
rect 82136 1244 84016 1272
rect 82136 1232 82142 1244
rect 84010 1232 84016 1244
rect 84068 1232 84074 1284
rect 84470 1232 84476 1284
rect 84528 1272 84534 1284
rect 86402 1272 86408 1284
rect 84528 1244 86408 1272
rect 84528 1232 84534 1244
rect 86402 1232 86408 1244
rect 86460 1232 86466 1284
rect 90358 1232 90364 1284
rect 90416 1272 90422 1284
rect 92198 1272 92204 1284
rect 90416 1244 92204 1272
rect 90416 1232 90422 1244
rect 92198 1232 92204 1244
rect 92256 1232 92262 1284
rect 92750 1232 92756 1284
rect 92808 1272 92814 1284
rect 94498 1272 94504 1284
rect 92808 1244 94504 1272
rect 92808 1232 92814 1244
rect 94498 1232 94504 1244
rect 94556 1232 94562 1284
rect 98638 1232 98644 1284
rect 98696 1272 98702 1284
rect 100294 1272 100300 1284
rect 98696 1244 100300 1272
rect 98696 1232 98702 1244
rect 100294 1232 100300 1244
rect 100352 1232 100358 1284
rect 102226 1232 102232 1284
rect 102284 1272 102290 1284
rect 103790 1272 103796 1284
rect 102284 1244 103796 1272
rect 102284 1232 102290 1244
rect 103790 1232 103796 1244
rect 103848 1232 103854 1284
rect 108114 1232 108120 1284
rect 108172 1272 108178 1284
rect 109586 1272 109592 1284
rect 108172 1244 109592 1272
rect 108172 1232 108178 1244
rect 109586 1232 109592 1244
rect 109644 1232 109650 1284
rect 110506 1232 110512 1284
rect 110564 1272 110570 1284
rect 111886 1272 111892 1284
rect 110564 1244 111892 1272
rect 110564 1232 110570 1244
rect 111886 1232 111892 1244
rect 111944 1232 111950 1284
rect 115198 1232 115204 1284
rect 115256 1272 115262 1284
rect 116578 1272 116584 1284
rect 115256 1244 116584 1272
rect 115256 1232 115262 1244
rect 116578 1232 116584 1244
rect 116636 1232 116642 1284
rect 117590 1232 117596 1284
rect 117648 1272 117654 1284
rect 118878 1272 118884 1284
rect 117648 1244 118884 1272
rect 117648 1232 117654 1244
rect 118878 1232 118884 1244
rect 118936 1232 118942 1284
rect 122282 1232 122288 1284
rect 122340 1272 122346 1284
rect 123478 1272 123484 1284
rect 122340 1244 123484 1272
rect 122340 1232 122346 1244
rect 123478 1232 123484 1244
rect 123536 1232 123542 1284
rect 124674 1232 124680 1284
rect 124732 1272 124738 1284
rect 125778 1272 125784 1284
rect 124732 1244 125784 1272
rect 124732 1232 124738 1244
rect 125778 1232 125784 1244
rect 125836 1232 125842 1284
rect 128170 1232 128176 1284
rect 128228 1272 128234 1284
rect 129274 1272 129280 1284
rect 128228 1244 129280 1272
rect 128228 1232 128234 1244
rect 129274 1232 129280 1244
rect 129332 1232 129338 1284
rect 136450 1232 136456 1284
rect 136508 1272 136514 1284
rect 137370 1272 137376 1284
rect 136508 1244 137376 1272
rect 136508 1232 136514 1244
rect 137370 1232 137376 1244
rect 137428 1232 137434 1284
rect 138842 1232 138848 1284
rect 138900 1272 138906 1284
rect 139762 1272 139768 1284
rect 138900 1244 139768 1272
rect 138900 1232 138906 1244
rect 139762 1232 139768 1244
rect 139820 1232 139826 1284
rect 140038 1232 140044 1284
rect 140096 1272 140102 1284
rect 140866 1272 140872 1284
rect 140096 1244 140872 1272
rect 140096 1232 140102 1244
rect 140866 1232 140872 1244
rect 140924 1232 140930 1284
rect 281350 1232 281356 1284
rect 281408 1272 281414 1284
rect 283098 1272 283104 1284
rect 281408 1244 283104 1272
rect 281408 1232 281414 1244
rect 283098 1232 283104 1244
rect 283156 1232 283162 1284
rect 289446 1232 289452 1284
rect 289504 1272 289510 1284
rect 291378 1272 291384 1284
rect 289504 1244 291384 1272
rect 289504 1232 289510 1244
rect 291378 1232 291384 1244
rect 291436 1232 291442 1284
rect 296438 1232 296444 1284
rect 296496 1272 296502 1284
rect 298462 1272 298468 1284
rect 296496 1244 298468 1272
rect 296496 1232 296502 1244
rect 298462 1232 298468 1244
rect 298520 1232 298526 1284
rect 303338 1232 303344 1284
rect 303396 1272 303402 1284
rect 305546 1272 305552 1284
rect 303396 1244 305552 1272
rect 303396 1232 303402 1244
rect 305546 1232 305552 1244
rect 305604 1232 305610 1284
rect 312538 1232 312544 1284
rect 312596 1272 312602 1284
rect 315022 1272 315028 1284
rect 312596 1244 315028 1272
rect 312596 1232 312602 1244
rect 315022 1232 315028 1244
rect 315080 1232 315086 1284
rect 318426 1232 318432 1284
rect 318484 1272 318490 1284
rect 320910 1272 320916 1284
rect 318484 1244 320916 1272
rect 318484 1232 318490 1244
rect 320910 1232 320916 1244
rect 320968 1232 320974 1284
rect 330018 1232 330024 1284
rect 330076 1272 330082 1284
rect 332686 1272 332692 1284
rect 330076 1244 332692 1272
rect 330076 1232 330082 1244
rect 332686 1232 332692 1244
rect 332744 1232 332750 1284
rect 334710 1232 334716 1284
rect 334768 1272 334774 1284
rect 337470 1272 337476 1284
rect 334768 1244 337476 1272
rect 334768 1232 334774 1244
rect 337470 1232 337476 1244
rect 337528 1232 337534 1284
rect 340506 1232 340512 1284
rect 340564 1272 340570 1284
rect 343358 1272 343364 1284
rect 340564 1244 343364 1272
rect 340564 1232 340570 1244
rect 343358 1232 343364 1244
rect 343416 1232 343422 1284
rect 344002 1232 344008 1284
rect 344060 1272 344066 1284
rect 346946 1272 346952 1284
rect 344060 1244 346952 1272
rect 344060 1232 344066 1244
rect 346946 1232 346952 1244
rect 347004 1232 347010 1284
rect 348602 1232 348608 1284
rect 348660 1272 348666 1284
rect 351638 1272 351644 1284
rect 348660 1244 351644 1272
rect 348660 1232 348666 1244
rect 351638 1232 351644 1244
rect 351696 1232 351702 1284
rect 352098 1232 352104 1284
rect 352156 1272 352162 1284
rect 355226 1272 355232 1284
rect 352156 1244 355232 1272
rect 352156 1232 352162 1244
rect 355226 1232 355232 1244
rect 355284 1232 355290 1284
rect 355594 1232 355600 1284
rect 355652 1272 355658 1284
rect 358722 1272 358728 1284
rect 355652 1244 358728 1272
rect 355652 1232 355658 1244
rect 358722 1232 358728 1244
rect 358780 1232 358786 1284
rect 359090 1232 359096 1284
rect 359148 1272 359154 1284
rect 362310 1272 362316 1284
rect 359148 1244 362316 1272
rect 359148 1232 359154 1244
rect 362310 1232 362316 1244
rect 362368 1232 362374 1284
rect 363690 1232 363696 1284
rect 363748 1272 363754 1284
rect 367002 1272 367008 1284
rect 363748 1244 367008 1272
rect 363748 1232 363754 1244
rect 367002 1232 367008 1244
rect 367060 1232 367066 1284
rect 372982 1232 372988 1284
rect 373040 1272 373046 1284
rect 376478 1272 376484 1284
rect 373040 1244 376484 1272
rect 373040 1232 373046 1244
rect 376478 1232 376484 1244
rect 376536 1232 376542 1284
rect 377582 1232 377588 1284
rect 377640 1272 377646 1284
rect 381170 1272 381176 1284
rect 377640 1244 381176 1272
rect 377640 1232 377646 1244
rect 381170 1232 381176 1244
rect 381228 1232 381234 1284
rect 388070 1232 388076 1284
rect 388128 1272 388134 1284
rect 391842 1272 391848 1284
rect 388128 1244 391848 1272
rect 388128 1232 388134 1244
rect 391842 1232 391848 1244
rect 391900 1232 391906 1284
rect 393866 1232 393872 1284
rect 393924 1272 393930 1284
rect 397730 1272 397736 1284
rect 393924 1244 397736 1272
rect 393924 1232 393930 1244
rect 397730 1232 397736 1244
rect 397788 1232 397794 1284
rect 403158 1232 403164 1284
rect 403216 1272 403222 1284
rect 407206 1272 407212 1284
rect 403216 1244 407212 1272
rect 403216 1232 403222 1244
rect 407206 1232 407212 1244
rect 407264 1232 407270 1284
rect 410058 1232 410064 1284
rect 410116 1272 410122 1284
rect 414290 1272 414296 1284
rect 410116 1244 414296 1272
rect 410116 1232 410122 1244
rect 414290 1232 414296 1244
rect 414348 1232 414354 1284
rect 418246 1232 418252 1284
rect 418304 1272 418310 1284
rect 422570 1272 422576 1284
rect 418304 1244 422576 1272
rect 418304 1232 418310 1244
rect 422570 1232 422576 1244
rect 422628 1232 422634 1284
rect 426342 1232 426348 1284
rect 426400 1272 426406 1284
rect 430850 1272 430856 1284
rect 426400 1244 430856 1272
rect 426400 1232 426406 1244
rect 430850 1232 430856 1244
rect 430908 1232 430914 1284
rect 435634 1232 435640 1284
rect 435692 1272 435698 1284
rect 439958 1272 439964 1284
rect 435692 1244 439964 1272
rect 435692 1232 435698 1244
rect 439958 1232 439964 1244
rect 440016 1232 440022 1284
rect 443730 1232 443736 1284
rect 443788 1272 443794 1284
rect 448238 1272 448244 1284
rect 443788 1244 448244 1272
rect 443788 1232 443794 1244
rect 448238 1232 448244 1244
rect 448296 1232 448302 1284
rect 450722 1232 450728 1284
rect 450780 1272 450786 1284
rect 455690 1272 455696 1284
rect 450780 1244 455696 1272
rect 450780 1232 450786 1244
rect 455690 1232 455696 1244
rect 455748 1232 455754 1284
rect 456518 1232 456524 1284
rect 456576 1272 456582 1284
rect 461578 1272 461584 1284
rect 456576 1244 461584 1272
rect 456576 1232 456582 1244
rect 461578 1232 461584 1244
rect 461636 1232 461642 1284
rect 462222 1232 462228 1284
rect 462280 1272 462286 1284
rect 467466 1272 467472 1284
rect 462280 1244 467472 1272
rect 462280 1232 462286 1244
rect 467466 1232 467472 1244
rect 467524 1232 467530 1284
rect 471606 1232 471612 1284
rect 471664 1272 471670 1284
rect 476574 1272 476580 1284
rect 471664 1244 476580 1272
rect 471664 1232 471670 1244
rect 476574 1232 476580 1244
rect 476632 1232 476638 1284
rect 480898 1232 480904 1284
rect 480956 1272 480962 1284
rect 486418 1272 486424 1284
rect 480956 1244 486424 1272
rect 480956 1232 480962 1244
rect 486418 1232 486424 1244
rect 486476 1232 486482 1284
rect 492490 1232 492496 1284
rect 492548 1272 492554 1284
rect 498194 1272 498200 1284
rect 492548 1244 498200 1272
rect 492548 1232 492554 1244
rect 498194 1232 498200 1244
rect 498252 1232 498258 1284
rect 498286 1232 498292 1284
rect 498344 1272 498350 1284
rect 503806 1272 503812 1284
rect 498344 1244 503812 1272
rect 498344 1232 498350 1244
rect 503806 1232 503812 1244
rect 503864 1232 503870 1284
rect 509878 1232 509884 1284
rect 509936 1272 509942 1284
rect 515582 1272 515588 1284
rect 509936 1244 515588 1272
rect 509936 1232 509942 1244
rect 515582 1232 515588 1244
rect 515640 1232 515646 1284
rect 517974 1232 517980 1284
rect 518032 1272 518038 1284
rect 523862 1272 523868 1284
rect 518032 1244 523868 1272
rect 518032 1232 518038 1244
rect 523862 1232 523868 1244
rect 523920 1232 523926 1284
rect 527266 1232 527272 1284
rect 527324 1272 527330 1284
rect 533706 1272 533712 1284
rect 527324 1244 533712 1272
rect 527324 1232 527330 1244
rect 533706 1232 533712 1244
rect 533764 1232 533770 1284
rect 537662 1232 537668 1284
rect 537720 1272 537726 1284
rect 544378 1272 544384 1284
rect 537720 1244 544384 1272
rect 537720 1232 537726 1244
rect 544378 1232 544384 1244
rect 544436 1232 544442 1284
rect 549346 1232 549352 1284
rect 549404 1272 549410 1284
rect 556154 1272 556160 1284
rect 549404 1244 556160 1272
rect 549404 1232 549410 1244
rect 556154 1232 556160 1244
rect 556212 1232 556218 1284
rect 563238 1232 563244 1284
rect 563296 1272 563302 1284
rect 570322 1272 570328 1284
rect 563296 1244 570328 1272
rect 563296 1232 563302 1244
rect 570322 1232 570328 1244
rect 570380 1232 570386 1284
rect 571260 1272 571288 1312
rect 572530 1300 572536 1352
rect 572588 1340 572594 1352
rect 579430 1340 579436 1352
rect 572588 1312 579436 1340
rect 572588 1300 572594 1312
rect 579430 1300 579436 1312
rect 579488 1300 579494 1352
rect 573542 1272 573548 1284
rect 571260 1244 573548 1272
rect 573542 1232 573548 1244
rect 573600 1232 573606 1284
rect 576118 1232 576124 1284
rect 576176 1272 576182 1284
rect 583386 1272 583392 1284
rect 576176 1244 583392 1272
rect 576176 1232 576182 1244
rect 583386 1232 583392 1244
rect 583444 1232 583450 1284
rect 99834 1164 99840 1216
rect 99892 1204 99898 1216
rect 101490 1204 101496 1216
rect 99892 1176 101496 1204
rect 99892 1164 99898 1176
rect 101490 1164 101496 1176
rect 101548 1164 101554 1216
rect 114002 1164 114008 1216
rect 114060 1204 114066 1216
rect 115382 1204 115388 1216
rect 114060 1176 115388 1204
rect 114060 1164 114066 1176
rect 115382 1164 115388 1176
rect 115440 1164 115446 1216
rect 311526 1164 311532 1216
rect 311584 1204 311590 1216
rect 313826 1204 313832 1216
rect 311584 1176 313832 1204
rect 311584 1164 311590 1176
rect 313826 1164 313832 1176
rect 313884 1164 313890 1216
rect 319622 1164 319628 1216
rect 319680 1204 319686 1216
rect 322106 1204 322112 1216
rect 319680 1176 322112 1204
rect 319680 1164 319686 1176
rect 322106 1164 322112 1176
rect 322164 1164 322170 1216
rect 327718 1164 327724 1216
rect 327776 1204 327782 1216
rect 330386 1204 330392 1216
rect 327776 1176 330392 1204
rect 327776 1164 327782 1176
rect 330386 1164 330392 1176
rect 330444 1164 330450 1216
rect 331122 1164 331128 1216
rect 331180 1204 331186 1216
rect 333882 1204 333888 1216
rect 331180 1176 333888 1204
rect 331180 1164 331186 1176
rect 333882 1164 333888 1176
rect 333940 1164 333946 1216
rect 337010 1164 337016 1216
rect 337068 1204 337074 1216
rect 339862 1204 339868 1216
rect 337068 1176 339868 1204
rect 337068 1164 337074 1176
rect 339862 1164 339868 1176
rect 339920 1164 339926 1216
rect 341702 1164 341708 1216
rect 341760 1204 341766 1216
rect 344554 1204 344560 1216
rect 341760 1176 344560 1204
rect 341760 1164 341766 1176
rect 344554 1164 344560 1176
rect 344612 1164 344618 1216
rect 357894 1164 357900 1216
rect 357952 1204 357958 1216
rect 361114 1204 361120 1216
rect 357952 1176 361120 1204
rect 357952 1164 357958 1176
rect 361114 1164 361120 1176
rect 361172 1164 361178 1216
rect 364886 1164 364892 1216
rect 364944 1204 364950 1216
rect 368198 1204 368204 1216
rect 364944 1176 368204 1204
rect 364944 1164 364950 1176
rect 368198 1164 368204 1176
rect 368256 1164 368262 1216
rect 375282 1164 375288 1216
rect 375340 1204 375346 1216
rect 378870 1204 378876 1216
rect 375340 1176 378876 1204
rect 375340 1164 375346 1176
rect 378870 1164 378876 1176
rect 378928 1164 378934 1216
rect 381078 1164 381084 1216
rect 381136 1204 381142 1216
rect 384758 1204 384764 1216
rect 381136 1176 384764 1204
rect 381136 1164 381142 1176
rect 384758 1164 384764 1176
rect 384816 1164 384822 1216
rect 390370 1164 390376 1216
rect 390428 1204 390434 1216
rect 394234 1204 394240 1216
rect 390428 1176 394240 1204
rect 390428 1164 390434 1176
rect 394234 1164 394240 1176
rect 394292 1164 394298 1216
rect 396166 1164 396172 1216
rect 396224 1204 396230 1216
rect 400122 1204 400128 1216
rect 396224 1176 400128 1204
rect 396224 1164 396230 1176
rect 400122 1164 400128 1176
rect 400180 1164 400186 1216
rect 400858 1164 400864 1216
rect 400916 1204 400922 1216
rect 404814 1204 404820 1216
rect 400916 1176 404820 1204
rect 400916 1164 400922 1176
rect 404814 1164 404820 1176
rect 404872 1164 404878 1216
rect 407758 1164 407764 1216
rect 407816 1204 407822 1216
rect 411898 1204 411904 1216
rect 407816 1176 411904 1204
rect 407816 1164 407822 1176
rect 411898 1164 411904 1176
rect 411956 1164 411962 1216
rect 420546 1164 420552 1216
rect 420604 1204 420610 1216
rect 424962 1204 424968 1216
rect 420604 1176 424968 1204
rect 420604 1164 420610 1176
rect 424962 1164 424968 1176
rect 425020 1164 425026 1216
rect 425146 1164 425152 1216
rect 425204 1204 425210 1216
rect 429654 1204 429660 1216
rect 425204 1176 429660 1204
rect 425204 1164 425210 1176
rect 429654 1164 429660 1176
rect 429712 1164 429718 1216
rect 441430 1164 441436 1216
rect 441488 1204 441494 1216
rect 445846 1204 445852 1216
rect 441488 1176 445852 1204
rect 441488 1164 441494 1176
rect 445846 1164 445852 1176
rect 445904 1164 445910 1216
rect 447226 1164 447232 1216
rect 447284 1204 447290 1216
rect 452102 1204 452108 1216
rect 447284 1176 452108 1204
rect 447284 1164 447290 1176
rect 452102 1164 452108 1176
rect 452160 1164 452166 1216
rect 454218 1164 454224 1216
rect 454276 1204 454282 1216
rect 459186 1204 459192 1216
rect 454276 1176 459192 1204
rect 454276 1164 454282 1176
rect 459186 1164 459192 1176
rect 459244 1164 459250 1216
rect 460014 1164 460020 1216
rect 460072 1204 460078 1216
rect 464798 1204 464804 1216
rect 460072 1176 464804 1204
rect 460072 1164 460078 1176
rect 464798 1164 464804 1176
rect 464856 1164 464862 1216
rect 470410 1164 470416 1216
rect 470468 1204 470474 1216
rect 475746 1204 475752 1216
rect 470468 1176 475752 1204
rect 470468 1164 470474 1176
rect 475746 1164 475752 1176
rect 475804 1164 475810 1216
rect 477402 1164 477408 1216
rect 477460 1204 477466 1216
rect 482462 1204 482468 1216
rect 477460 1176 482468 1204
rect 477460 1164 477466 1176
rect 482462 1164 482468 1176
rect 482520 1164 482526 1216
rect 483198 1164 483204 1216
rect 483256 1204 483262 1216
rect 488810 1204 488816 1216
rect 483256 1176 488816 1204
rect 483256 1164 483262 1176
rect 488810 1164 488816 1176
rect 488868 1164 488874 1216
rect 490098 1164 490104 1216
rect 490156 1204 490162 1216
rect 495526 1204 495532 1216
rect 490156 1176 495532 1204
rect 490156 1164 490162 1176
rect 495526 1164 495532 1176
rect 495584 1164 495590 1216
rect 505186 1164 505192 1216
rect 505244 1204 505250 1216
rect 511258 1204 511264 1216
rect 505244 1176 511264 1204
rect 505244 1164 505250 1176
rect 511258 1164 511264 1176
rect 511316 1164 511322 1216
rect 514478 1164 514484 1216
rect 514536 1204 514542 1216
rect 520366 1204 520372 1216
rect 514536 1176 520372 1204
rect 514536 1164 514542 1176
rect 520366 1164 520372 1176
rect 520424 1164 520430 1216
rect 521470 1164 521476 1216
rect 521528 1204 521534 1216
rect 527818 1204 527824 1216
rect 521528 1176 527824 1204
rect 521528 1164 521534 1176
rect 527818 1164 527824 1176
rect 527876 1164 527882 1216
rect 528462 1164 528468 1216
rect 528520 1204 528526 1216
rect 534534 1204 534540 1216
rect 528520 1176 534540 1204
rect 528520 1164 528526 1176
rect 534534 1164 534540 1176
rect 534592 1164 534598 1216
rect 542262 1164 542268 1216
rect 542320 1204 542326 1216
rect 548702 1204 548708 1216
rect 542320 1176 548708 1204
rect 542320 1164 542326 1176
rect 548702 1164 548708 1176
rect 548760 1164 548766 1216
rect 556246 1164 556252 1216
rect 556304 1204 556310 1216
rect 563146 1204 563152 1216
rect 556304 1176 563152 1204
rect 556304 1164 556310 1176
rect 563146 1164 563152 1176
rect 563204 1164 563210 1216
rect 569034 1164 569040 1216
rect 569092 1204 569098 1216
rect 575934 1204 575940 1216
rect 569092 1176 575940 1204
rect 569092 1164 569098 1176
rect 575934 1164 575940 1176
rect 575992 1164 575998 1216
rect 5626 1096 5632 1148
rect 5684 1136 5690 1148
rect 8662 1136 8668 1148
rect 5684 1108 8668 1136
rect 5684 1096 5690 1108
rect 8662 1096 8668 1108
rect 8720 1096 8726 1148
rect 111610 1096 111616 1148
rect 111668 1136 111674 1148
rect 113082 1136 113088 1148
rect 111668 1108 113088 1136
rect 111668 1096 111674 1108
rect 113082 1096 113088 1108
rect 113140 1096 113146 1148
rect 123478 1096 123484 1148
rect 123536 1136 123542 1148
rect 124766 1136 124772 1148
rect 123536 1108 124772 1136
rect 123536 1096 123542 1108
rect 124766 1096 124772 1108
rect 124824 1096 124830 1148
rect 320818 1096 320824 1148
rect 320876 1136 320882 1148
rect 323302 1136 323308 1148
rect 320876 1108 323308 1136
rect 320876 1096 320882 1108
rect 323302 1096 323308 1108
rect 323360 1096 323366 1148
rect 360102 1096 360108 1148
rect 360160 1136 360166 1148
rect 363506 1136 363512 1148
rect 360160 1108 363512 1136
rect 360160 1096 360166 1108
rect 363506 1096 363512 1108
rect 363564 1096 363570 1148
rect 382182 1096 382188 1148
rect 382240 1136 382246 1148
rect 385954 1136 385960 1148
rect 382240 1108 385960 1136
rect 382240 1096 382246 1108
rect 385954 1096 385960 1108
rect 386012 1096 386018 1148
rect 389266 1096 389272 1148
rect 389324 1136 389330 1148
rect 393038 1136 393044 1148
rect 389324 1108 393044 1136
rect 389324 1096 389330 1108
rect 393038 1096 393044 1108
rect 393096 1096 393102 1148
rect 398466 1096 398472 1148
rect 398524 1136 398530 1148
rect 402514 1136 402520 1148
rect 398524 1108 402520 1136
rect 398524 1096 398530 1108
rect 402514 1096 402520 1108
rect 402572 1096 402578 1148
rect 404262 1096 404268 1148
rect 404320 1136 404326 1148
rect 408402 1136 408408 1148
rect 404320 1108 408408 1136
rect 404320 1096 404326 1108
rect 408402 1096 408408 1108
rect 408460 1096 408466 1148
rect 408954 1096 408960 1148
rect 409012 1136 409018 1148
rect 413094 1136 413100 1148
rect 409012 1108 413100 1136
rect 409012 1096 409018 1108
rect 413094 1096 413100 1108
rect 413152 1096 413158 1148
rect 415946 1096 415952 1148
rect 416004 1136 416010 1148
rect 420178 1136 420184 1148
rect 416004 1108 420184 1136
rect 416004 1096 416010 1108
rect 420178 1096 420184 1108
rect 420236 1096 420242 1148
rect 429838 1096 429844 1148
rect 429896 1136 429902 1148
rect 434438 1136 434444 1148
rect 429896 1108 434444 1136
rect 429896 1096 429902 1108
rect 434438 1096 434444 1108
rect 434496 1096 434502 1148
rect 436738 1096 436744 1148
rect 436796 1136 436802 1148
rect 441522 1136 441528 1148
rect 436796 1108 441528 1136
rect 436796 1096 436802 1108
rect 441522 1096 441528 1108
rect 441580 1096 441586 1148
rect 446030 1096 446036 1148
rect 446088 1136 446094 1148
rect 450906 1136 450912 1148
rect 446088 1108 450912 1136
rect 446088 1096 446094 1108
rect 450906 1096 450912 1108
rect 450964 1096 450970 1148
rect 457622 1096 457628 1148
rect 457680 1136 457686 1148
rect 462406 1136 462412 1148
rect 457680 1108 462412 1136
rect 457680 1096 457686 1108
rect 462406 1096 462412 1108
rect 462464 1096 462470 1148
rect 464614 1096 464620 1148
rect 464672 1136 464678 1148
rect 469858 1136 469864 1148
rect 464672 1108 469864 1136
rect 464672 1096 464678 1108
rect 469858 1096 469864 1108
rect 469916 1096 469922 1148
rect 472710 1096 472716 1148
rect 472768 1136 472774 1148
rect 478138 1136 478144 1148
rect 472768 1108 478144 1136
rect 472768 1096 472774 1108
rect 478138 1096 478144 1108
rect 478196 1096 478202 1148
rect 486694 1096 486700 1148
rect 486752 1136 486758 1148
rect 492306 1136 492312 1148
rect 486752 1108 492312 1136
rect 486752 1096 486758 1108
rect 492306 1096 492312 1108
rect 492364 1096 492370 1148
rect 500586 1096 500592 1148
rect 500644 1136 500650 1148
rect 506474 1136 506480 1148
rect 500644 1108 506480 1136
rect 500644 1096 500650 1108
rect 506474 1096 506480 1108
rect 506532 1096 506538 1148
rect 510982 1096 510988 1148
rect 511040 1136 511046 1148
rect 517146 1136 517152 1148
rect 511040 1108 517152 1136
rect 511040 1096 511046 1108
rect 517146 1096 517152 1108
rect 517204 1096 517210 1148
rect 522666 1096 522672 1148
rect 522724 1136 522730 1148
rect 528646 1136 528652 1148
rect 522724 1108 528652 1136
rect 522724 1096 522730 1108
rect 528646 1096 528652 1108
rect 528704 1096 528710 1148
rect 530762 1096 530768 1148
rect 530820 1136 530826 1148
rect 537202 1136 537208 1148
rect 530820 1108 537208 1136
rect 530820 1096 530826 1108
rect 537202 1096 537208 1108
rect 537260 1096 537266 1148
rect 543458 1096 543464 1148
rect 543516 1136 543522 1148
rect 550266 1136 550272 1148
rect 543516 1108 550272 1136
rect 543516 1096 543522 1108
rect 550266 1096 550272 1108
rect 550324 1096 550330 1148
rect 550450 1096 550456 1148
rect 550508 1136 550514 1148
rect 556982 1136 556988 1148
rect 550508 1108 556988 1136
rect 550508 1096 550514 1108
rect 556982 1096 556988 1108
rect 557040 1096 557046 1148
rect 558546 1096 558552 1148
rect 558604 1136 558610 1148
rect 565262 1136 565268 1148
rect 558604 1108 565268 1136
rect 558604 1096 558610 1108
rect 565262 1096 565268 1108
rect 565320 1096 565326 1148
rect 567838 1096 567844 1148
rect 567896 1136 567902 1148
rect 575106 1136 575112 1148
rect 567896 1108 575112 1136
rect 567896 1096 567902 1108
rect 575106 1096 575112 1108
rect 575164 1096 575170 1148
rect 378778 1028 378784 1080
rect 378836 1068 378842 1080
rect 382366 1068 382372 1080
rect 378836 1040 382372 1068
rect 378836 1028 378842 1040
rect 382366 1028 382372 1040
rect 382424 1028 382430 1080
rect 386874 1028 386880 1080
rect 386932 1068 386938 1080
rect 390646 1068 390652 1080
rect 386932 1040 390652 1068
rect 386932 1028 386938 1040
rect 390646 1028 390652 1040
rect 390704 1028 390710 1080
rect 417050 1028 417056 1080
rect 417108 1068 417114 1080
rect 421374 1068 421380 1080
rect 417108 1040 421380 1068
rect 417108 1028 417114 1040
rect 421374 1028 421380 1040
rect 421432 1028 421438 1080
rect 428642 1028 428648 1080
rect 428700 1068 428706 1080
rect 433242 1068 433248 1080
rect 428700 1040 433248 1068
rect 428700 1028 428706 1040
rect 433242 1028 433248 1040
rect 433300 1028 433306 1080
rect 437934 1028 437940 1080
rect 437992 1068 437998 1080
rect 442626 1068 442632 1080
rect 437992 1040 442632 1068
rect 437992 1028 437998 1040
rect 442626 1028 442632 1040
rect 442684 1028 442690 1080
rect 455322 1028 455328 1080
rect 455380 1068 455386 1080
rect 460014 1068 460020 1080
rect 455380 1040 460020 1068
rect 455380 1028 455386 1040
rect 460014 1028 460020 1040
rect 460072 1028 460078 1080
rect 465810 1028 465816 1080
rect 465868 1068 465874 1080
rect 470686 1068 470692 1080
rect 465868 1040 470692 1068
rect 465868 1028 465874 1040
rect 470686 1028 470692 1040
rect 470744 1028 470750 1080
rect 473906 1028 473912 1080
rect 473964 1068 473970 1080
rect 478966 1068 478972 1080
rect 473964 1040 478972 1068
rect 473964 1028 473970 1040
rect 478966 1028 478972 1040
rect 479024 1028 479030 1080
rect 482002 1028 482008 1080
rect 482060 1068 482066 1080
rect 487246 1068 487252 1080
rect 482060 1040 487252 1068
rect 482060 1028 482066 1040
rect 487246 1028 487252 1040
rect 487304 1028 487310 1080
rect 491202 1028 491208 1080
rect 491260 1068 491266 1080
rect 497090 1068 497096 1080
rect 491260 1040 497096 1068
rect 491260 1028 491266 1040
rect 497090 1028 497096 1040
rect 497148 1028 497154 1080
rect 499390 1028 499396 1080
rect 499448 1068 499454 1080
rect 505370 1068 505376 1080
rect 499448 1040 505376 1068
rect 499448 1028 499454 1040
rect 505370 1028 505376 1040
rect 505428 1028 505434 1080
rect 508682 1028 508688 1080
rect 508740 1068 508746 1080
rect 514754 1068 514760 1080
rect 508740 1040 514760 1068
rect 508740 1028 508746 1040
rect 514754 1028 514760 1040
rect 514812 1028 514818 1080
rect 519170 1028 519176 1080
rect 519228 1068 519234 1080
rect 525426 1068 525432 1080
rect 519228 1040 525432 1068
rect 519228 1028 519234 1040
rect 525426 1028 525432 1040
rect 525484 1028 525490 1080
rect 531866 1028 531872 1080
rect 531924 1068 531930 1080
rect 538214 1068 538220 1080
rect 531924 1040 538220 1068
rect 531924 1028 531930 1040
rect 538214 1028 538220 1040
rect 538272 1028 538278 1080
rect 538858 1028 538864 1080
rect 538916 1068 538922 1080
rect 545482 1068 545488 1080
rect 538916 1040 545488 1068
rect 538916 1028 538922 1040
rect 545482 1028 545488 1040
rect 545540 1028 545546 1080
rect 546954 1028 546960 1080
rect 547012 1068 547018 1080
rect 553762 1068 553768 1080
rect 547012 1040 553768 1068
rect 547012 1028 547018 1040
rect 553762 1028 553768 1040
rect 553820 1028 553826 1080
rect 560938 1028 560944 1080
rect 560996 1068 561002 1080
rect 567654 1068 567660 1080
rect 560996 1040 567660 1068
rect 560996 1028 561002 1040
rect 567654 1028 567660 1040
rect 567712 1028 567718 1080
rect 571242 1028 571248 1080
rect 571300 1068 571306 1080
rect 578602 1068 578608 1080
rect 571300 1040 578608 1068
rect 571300 1028 571306 1040
rect 578602 1028 578608 1040
rect 578660 1028 578666 1080
rect 326614 960 326620 1012
rect 326672 1000 326678 1012
rect 329190 1000 329196 1012
rect 326672 972 329196 1000
rect 326672 960 326678 972
rect 329190 960 329196 972
rect 329248 960 329254 1012
rect 374178 960 374184 1012
rect 374236 1000 374242 1012
rect 377674 1000 377680 1012
rect 374236 972 377680 1000
rect 374236 960 374242 972
rect 377674 960 377680 972
rect 377732 960 377738 1012
rect 379882 960 379888 1012
rect 379940 1000 379946 1012
rect 383562 1000 383568 1012
rect 379940 972 383568 1000
rect 379940 960 379946 972
rect 383562 960 383568 972
rect 383620 960 383626 1012
rect 414750 960 414756 1012
rect 414808 1000 414814 1012
rect 418982 1000 418988 1012
rect 414808 972 418988 1000
rect 414808 960 414814 972
rect 418982 960 418988 972
rect 419040 960 419046 1012
rect 424042 960 424048 1012
rect 424100 1000 424106 1012
rect 428458 1000 428464 1012
rect 424100 972 428464 1000
rect 424100 960 424106 972
rect 428458 960 428464 972
rect 428516 960 428522 1012
rect 432138 960 432144 1012
rect 432196 1000 432202 1012
rect 436738 1000 436744 1012
rect 432196 972 436744 1000
rect 432196 960 432202 972
rect 436738 960 436744 972
rect 436796 960 436802 1012
rect 439130 960 439136 1012
rect 439188 1000 439194 1012
rect 443822 1000 443828 1012
rect 439188 972 443828 1000
rect 439188 960 439194 972
rect 443822 960 443828 972
rect 443880 960 443886 1012
rect 453022 960 453028 1012
rect 453080 1000 453086 1012
rect 458082 1000 458088 1012
rect 453080 972 458088 1000
rect 453080 960 453086 972
rect 458082 960 458088 972
rect 458140 960 458146 1012
rect 466914 960 466920 1012
rect 466972 1000 466978 1012
rect 472250 1000 472256 1012
rect 466972 972 472256 1000
rect 466972 960 466978 972
rect 472250 960 472256 972
rect 472308 960 472314 1012
rect 476206 960 476212 1012
rect 476264 1000 476270 1012
rect 481358 1000 481364 1012
rect 476264 972 481364 1000
rect 476264 960 476270 972
rect 481358 960 481364 972
rect 481416 960 481422 1012
rect 488994 960 489000 1012
rect 489052 1000 489058 1012
rect 494698 1000 494704 1012
rect 489052 972 494704 1000
rect 489052 960 489058 972
rect 494698 960 494704 972
rect 494756 960 494762 1012
rect 494790 960 494796 1012
rect 494848 1000 494854 1012
rect 500586 1000 500592 1012
rect 494848 972 500592 1000
rect 494848 960 494854 972
rect 500586 960 500592 972
rect 500644 960 500650 1012
rect 501782 960 501788 1012
rect 501840 1000 501846 1012
rect 507302 1000 507308 1012
rect 501840 972 507308 1000
rect 501840 960 501846 972
rect 507302 960 507308 972
rect 507360 960 507366 1012
rect 512178 960 512184 1012
rect 512236 1000 512242 1012
rect 517974 1000 517980 1012
rect 512236 972 517980 1000
rect 512236 960 512242 972
rect 517974 960 517980 972
rect 518032 960 518038 1012
rect 523770 960 523776 1012
rect 523828 1000 523834 1012
rect 529934 1000 529940 1012
rect 523828 972 529940 1000
rect 523828 960 523834 972
rect 529934 960 529940 972
rect 529992 960 529998 1012
rect 533062 960 533068 1012
rect 533120 1000 533126 1012
rect 539594 1000 539600 1012
rect 533120 972 539600 1000
rect 533120 960 533126 972
rect 539594 960 539600 972
rect 539652 960 539658 1012
rect 540054 960 540060 1012
rect 540112 1000 540118 1012
rect 546494 1000 546500 1012
rect 540112 972 546500 1000
rect 540112 960 540118 972
rect 546494 960 546500 972
rect 546552 960 546558 1012
rect 551646 960 551652 1012
rect 551704 1000 551710 1012
rect 558546 1000 558552 1012
rect 551704 972 558552 1000
rect 551704 960 551710 972
rect 558546 960 558552 972
rect 558604 960 558610 1012
rect 561950 960 561956 1012
rect 562008 1000 562014 1012
rect 568758 1000 568764 1012
rect 562008 972 568764 1000
rect 562008 960 562014 972
rect 568758 960 568764 972
rect 568816 960 568822 1012
rect 570138 960 570144 1012
rect 570196 1000 570202 1012
rect 577038 1000 577044 1012
rect 570196 972 577044 1000
rect 570196 960 570202 972
rect 577038 960 577044 972
rect 577096 960 577102 1012
rect 8754 892 8760 944
rect 8812 932 8818 944
rect 12158 932 12164 944
rect 8812 904 12164 932
rect 8812 892 8818 904
rect 12158 892 12164 904
rect 12216 892 12222 944
rect 121086 892 121092 944
rect 121144 932 121150 944
rect 122374 932 122380 944
rect 121144 904 122380 932
rect 121144 892 121150 904
rect 122374 892 122380 904
rect 122432 892 122438 944
rect 463418 892 463424 944
rect 463476 932 463482 944
rect 468294 932 468300 944
rect 463476 904 468300 932
rect 463476 892 463482 904
rect 468294 892 468300 904
rect 468352 892 468358 944
rect 479702 892 479708 944
rect 479760 932 479766 944
rect 484854 932 484860 944
rect 479760 904 484860 932
rect 479760 892 479766 904
rect 484854 892 484860 904
rect 484912 892 484918 944
rect 493594 892 493600 944
rect 493652 932 493658 944
rect 499390 932 499396 944
rect 493652 904 499396 932
rect 493652 892 493658 904
rect 499390 892 499396 904
rect 499448 892 499454 944
rect 502886 892 502892 944
rect 502944 932 502950 944
rect 508866 932 508872 944
rect 502944 904 508872 932
rect 502944 892 502950 904
rect 508866 892 508872 904
rect 508924 892 508930 944
rect 520182 892 520188 944
rect 520240 932 520246 944
rect 526254 932 526260 944
rect 520240 904 526260 932
rect 520240 892 520246 904
rect 526254 892 526260 904
rect 526312 892 526318 944
rect 529566 892 529572 944
rect 529624 932 529630 944
rect 536098 932 536104 944
rect 529624 904 536104 932
rect 529624 892 529630 904
rect 536098 892 536104 904
rect 536156 892 536162 944
rect 559650 892 559656 944
rect 559708 932 559714 944
rect 566826 932 566832 944
rect 559708 904 566832 932
rect 559708 892 559714 904
rect 566826 892 566832 904
rect 566884 892 566890 944
rect 347498 824 347504 876
rect 347556 864 347562 876
rect 350442 864 350448 876
rect 347556 836 350448 864
rect 347556 824 347562 836
rect 350442 824 350448 836
rect 350500 824 350506 876
rect 361390 824 361396 876
rect 361448 864 361454 876
rect 364610 864 364616 876
rect 361448 836 364616 864
rect 361448 824 361454 836
rect 364610 824 364616 836
rect 364668 824 364674 876
rect 368382 824 368388 876
rect 368440 864 368446 876
rect 371694 864 371700 876
rect 368440 836 371700 864
rect 368440 824 368446 836
rect 371694 824 371700 836
rect 371752 824 371758 876
rect 371786 824 371792 876
rect 371844 864 371850 876
rect 375282 864 375288 876
rect 371844 836 375288 864
rect 371844 824 371850 836
rect 375282 824 375288 836
rect 375340 824 375346 876
rect 384574 824 384580 876
rect 384632 864 384638 876
rect 388254 864 388260 876
rect 384632 836 388260 864
rect 384632 824 384638 836
rect 388254 824 388260 836
rect 388312 824 388318 876
rect 391566 824 391572 876
rect 391624 864 391630 876
rect 395338 864 395344 876
rect 391624 836 395344 864
rect 391624 824 391630 836
rect 395338 824 395344 836
rect 395396 824 395402 876
rect 397362 824 397368 876
rect 397420 864 397426 876
rect 401318 864 401324 876
rect 397420 836 401324 864
rect 397420 824 397426 836
rect 401318 824 401324 836
rect 401376 824 401382 876
rect 406654 824 406660 876
rect 406712 864 406718 876
rect 410794 864 410800 876
rect 406712 836 410800 864
rect 406712 824 406718 836
rect 410794 824 410800 836
rect 410852 824 410858 876
rect 419350 824 419356 876
rect 419408 864 419414 876
rect 423398 864 423404 876
rect 419408 836 423404 864
rect 419408 824 419414 836
rect 423398 824 423404 836
rect 423456 824 423462 876
rect 434346 824 434352 876
rect 434404 864 434410 876
rect 439130 864 439136 876
rect 434404 836 439136 864
rect 434404 824 434410 836
rect 439130 824 439136 836
rect 439188 824 439194 876
rect 444926 824 444932 876
rect 444984 864 444990 876
rect 449802 864 449808 876
rect 444984 836 449808 864
rect 444984 824 444990 836
rect 449802 824 449808 836
rect 449860 824 449866 876
rect 461118 824 461124 876
rect 461176 864 461182 876
rect 466270 864 466276 876
rect 461176 836 466276 864
rect 461176 824 461182 836
rect 466270 824 466276 836
rect 466328 824 466334 876
rect 484302 824 484308 876
rect 484360 864 484366 876
rect 489914 864 489920 876
rect 484360 836 489920 864
rect 484360 824 484366 836
rect 489914 824 489920 836
rect 489972 824 489978 876
rect 495986 824 495992 876
rect 496044 864 496050 876
rect 501782 864 501788 876
rect 496044 836 501788 864
rect 496044 824 496050 836
rect 501782 824 501788 836
rect 501840 824 501846 876
rect 552750 824 552756 876
rect 552808 864 552814 876
rect 559742 864 559748 876
rect 552808 836 559748 864
rect 552808 824 552814 836
rect 559742 824 559748 836
rect 559800 824 559806 876
rect 52546 688 52552 740
rect 52604 728 52610 740
rect 55030 728 55036 740
rect 52604 700 55036 728
rect 52604 688 52610 700
rect 55030 688 55036 700
rect 55088 688 55094 740
rect 59630 688 59636 740
rect 59688 728 59694 740
rect 61930 728 61936 740
rect 59688 700 61936 728
rect 59688 688 59694 700
rect 61930 688 61936 700
rect 61988 688 61994 740
rect 105722 688 105728 740
rect 105780 728 105786 740
rect 107286 728 107292 740
rect 105780 700 107292 728
rect 105780 688 105786 700
rect 107286 688 107292 700
rect 107344 688 107350 740
rect 274358 688 274364 740
rect 274416 728 274422 740
rect 276014 728 276020 740
rect 274416 700 276020 728
rect 274416 688 274422 700
rect 276014 688 276020 700
rect 276072 688 276078 740
rect 333514 688 333520 740
rect 333572 728 333578 740
rect 336274 728 336280 740
rect 333572 700 336280 728
rect 333572 688 333578 700
rect 336274 688 336280 700
rect 336332 688 336338 740
rect 338206 688 338212 740
rect 338264 728 338270 740
rect 340966 728 340972 740
rect 338264 700 340972 728
rect 338264 688 338270 700
rect 340966 688 340972 700
rect 341024 688 341030 740
rect 342806 688 342812 740
rect 342864 728 342870 740
rect 345750 728 345756 740
rect 342864 700 345756 728
rect 342864 688 342870 700
rect 345750 688 345756 700
rect 345808 688 345814 740
rect 346302 688 346308 740
rect 346360 728 346366 740
rect 349246 728 349252 740
rect 346360 700 349252 728
rect 346360 688 346366 700
rect 349246 688 349252 700
rect 349304 688 349310 740
rect 350902 688 350908 740
rect 350960 728 350966 740
rect 354030 728 354036 740
rect 350960 700 354036 728
rect 350960 688 350966 700
rect 354030 688 354036 700
rect 354088 688 354094 740
rect 365990 688 365996 740
rect 366048 728 366054 740
rect 369394 728 369400 740
rect 366048 700 369400 728
rect 366048 688 366054 700
rect 369394 688 369400 700
rect 369452 688 369458 740
rect 369486 688 369492 740
rect 369544 728 369550 740
rect 372890 728 372896 740
rect 369544 700 372896 728
rect 369544 688 369550 700
rect 372890 688 372896 700
rect 372948 688 372954 740
rect 451826 688 451832 740
rect 451884 728 451890 740
rect 456518 728 456524 740
rect 451884 700 456524 728
rect 451884 688 451890 700
rect 456518 688 456524 700
rect 456576 688 456582 740
rect 69106 552 69112 604
rect 69164 592 69170 604
rect 71314 592 71320 604
rect 69164 564 71320 592
rect 69164 552 69170 564
rect 71314 552 71320 564
rect 71372 552 71378 604
rect 290642 552 290648 604
rect 290700 592 290706 604
rect 292574 592 292580 604
rect 290700 564 292580 592
rect 290700 552 290706 564
rect 292574 552 292580 564
rect 292632 552 292638 604
rect 304534 552 304540 604
rect 304592 592 304598 604
rect 306742 592 306748 604
rect 304592 564 306748 592
rect 304592 552 304598 564
rect 306742 552 306748 564
rect 306800 552 306806 604
rect 324222 552 324228 604
rect 324280 592 324286 604
rect 326798 592 326804 604
rect 324280 564 326804 592
rect 324280 552 324286 564
rect 326798 552 326804 564
rect 326856 552 326862 604
rect 416682 552 416688 604
rect 416740 552 416746 604
rect 557534 552 557540 604
rect 557592 592 557598 604
rect 564434 592 564440 604
rect 557592 564 564440 592
rect 557592 552 557598 564
rect 564434 552 564440 564
rect 564492 552 564498 604
rect 412450 348 412456 400
rect 412508 388 412514 400
rect 416700 388 416728 552
rect 565446 416 565452 468
rect 565504 456 565510 468
rect 572898 456 572904 468
rect 565504 428 572904 456
rect 565504 416 565510 428
rect 572898 416 572904 428
rect 572956 416 572962 468
rect 412508 360 416728 388
rect 412508 348 412514 360
rect 401962 144 401968 196
rect 402020 184 402026 196
rect 406194 184 406200 196
rect 402020 156 406200 184
rect 402020 144 402026 156
rect 406194 144 406200 156
rect 406252 144 406258 196
rect 383378 76 383384 128
rect 383436 116 383442 128
rect 386782 116 386788 128
rect 383436 88 386788 116
rect 383436 76 383442 88
rect 386782 76 386788 88
rect 386840 76 386846 128
rect 421742 76 421748 128
rect 421800 116 421806 128
rect 425790 116 425796 128
rect 421800 88 425796 116
rect 421800 76 421806 88
rect 425790 76 425796 88
rect 425848 76 425854 128
rect 354398 8 354404 60
rect 354456 48 354462 60
rect 357342 48 357348 60
rect 354456 20 357348 48
rect 354456 8 354462 20
rect 357342 8 357348 20
rect 357400 8 357406 60
rect 392670 8 392676 60
rect 392728 48 392734 60
rect 396166 48 396172 60
rect 392728 20 396172 48
rect 392728 8 392734 20
rect 396166 8 396172 20
rect 396224 8 396230 60
rect 431034 8 431040 60
rect 431092 48 431098 60
rect 435174 48 435180 60
rect 431092 20 435180 48
rect 431092 8 431098 20
rect 435174 8 435180 20
rect 435232 8 435238 60
rect 469306 8 469312 60
rect 469364 48 469370 60
rect 474182 48 474188 60
rect 469364 20 474188 48
rect 469364 8 469370 20
rect 474182 8 474188 20
rect 474240 8 474246 60
rect 564250 8 564256 60
rect 564308 48 564314 60
rect 571334 48 571340 60
rect 564308 20 571340 48
rect 564308 8 564314 20
rect 571334 8 571340 20
rect 571392 8 571398 60
<< via1 >>
rect 3884 700748 3936 700800
rect 8116 700748 8168 700800
rect 348792 700544 348844 700596
rect 355876 700544 355928 700596
rect 105452 700272 105504 700324
rect 113916 700272 113968 700324
rect 170312 700272 170364 700324
rect 179880 700272 179932 700324
rect 218980 700272 219032 700324
rect 223856 700272 223908 700324
rect 235172 700272 235224 700324
rect 245844 700272 245896 700324
rect 283840 700272 283892 700324
rect 289820 700272 289872 700324
rect 300124 700272 300176 700324
rect 311900 700272 311952 700324
rect 364984 700272 365036 700324
rect 377864 700272 377916 700324
rect 429844 700272 429896 700324
rect 443828 700272 443880 700324
rect 478512 700272 478564 700324
rect 487804 700272 487856 700324
rect 494796 700272 494848 700324
rect 509792 700272 509844 700324
rect 527180 700272 527232 700324
rect 531780 700272 531832 700324
rect 543464 700272 543516 700324
rect 553768 700272 553820 700324
rect 559656 700272 559708 700324
rect 575756 700272 575808 700324
rect 24308 700204 24360 700256
rect 25964 700204 26016 700256
rect 40500 700204 40552 700256
rect 47952 700204 48004 700256
rect 70032 700204 70084 700256
rect 72976 700204 73028 700256
rect 89168 700204 89220 700256
rect 91928 700204 91980 700256
rect 135996 700204 136048 700256
rect 137836 700204 137888 700256
rect 154120 700204 154172 700256
rect 157892 700204 157944 700256
rect 201960 700204 202012 700256
rect 202788 700204 202840 700256
rect 397460 700204 397512 700256
rect 399852 700204 399904 700256
rect 413652 700204 413704 700256
rect 421840 700204 421892 700256
rect 462320 700204 462372 700256
rect 465816 700204 465868 700256
rect 332508 700068 332560 700120
rect 333888 700068 333940 700120
rect 578424 682456 578476 682508
rect 579988 682456 580040 682508
rect 20 423580 72 423632
rect 572 423580 624 423632
rect 578240 397468 578292 397520
rect 580264 397468 580316 397520
rect 578332 351024 578384 351076
rect 580264 351024 580316 351076
rect 578516 303696 578568 303748
rect 580264 303696 580316 303748
rect 578884 273164 578936 273216
rect 580816 273164 580868 273216
rect 578608 255280 578660 255332
rect 580264 255280 580316 255332
rect 578332 208360 578384 208412
rect 580264 208360 580316 208412
rect 578240 60664 578292 60716
rect 580816 60664 580868 60716
rect 11152 3884 11204 3936
rect 14508 3884 14560 3936
rect 14740 3884 14792 3936
rect 18004 3884 18056 3936
rect 20628 3884 20680 3936
rect 23800 3884 23852 3936
rect 24216 3884 24268 3936
rect 27296 3884 27348 3936
rect 27712 3884 27764 3936
rect 30700 3884 30752 3936
rect 32404 3884 32456 3936
rect 35392 3884 35444 3936
rect 38384 3884 38436 3936
rect 41188 3884 41240 3936
rect 43076 3884 43128 3936
rect 45788 3884 45840 3936
rect 46664 3884 46716 3936
rect 49284 3884 49336 3936
rect 50160 3884 50212 3936
rect 52780 3884 52832 3936
rect 56048 3884 56100 3936
rect 58576 3884 58628 3936
rect 72608 3884 72660 3936
rect 74860 3884 74912 3936
rect 247636 3884 247688 3936
rect 248604 3884 248656 3936
rect 285908 3884 285960 3936
rect 287796 3884 287848 3936
rect 1676 3816 1728 3868
rect 5216 3816 5268 3868
rect 13544 3816 13596 3868
rect 16808 3816 16860 3868
rect 19432 3816 19484 3868
rect 22604 3816 22656 3868
rect 23020 3816 23072 3868
rect 26100 3816 26152 3868
rect 26516 3816 26568 3868
rect 29596 3816 29648 3868
rect 30104 3816 30156 3868
rect 33092 3816 33144 3868
rect 33600 3816 33652 3868
rect 36588 3816 36640 3868
rect 37188 3816 37240 3868
rect 39992 3816 40044 3868
rect 41880 3816 41932 3868
rect 44684 3816 44736 3868
rect 45468 3816 45520 3868
rect 48180 3816 48232 3868
rect 48964 3816 49016 3868
rect 51584 3816 51636 3868
rect 53748 3816 53800 3868
rect 56276 3816 56328 3868
rect 57244 3816 57296 3868
rect 59772 3816 59824 3868
rect 71504 3816 71556 3868
rect 73664 3816 73716 3868
rect 78588 3816 78640 3868
rect 80656 3816 80708 3868
rect 80888 3816 80940 3868
rect 82956 3816 83008 3868
rect 87972 3816 88024 3868
rect 89948 3816 90000 3868
rect 96252 3816 96304 3868
rect 98044 3816 98096 3868
rect 244140 3816 244192 3868
rect 245200 3816 245252 3868
rect 256928 3816 256980 3868
rect 258264 3816 258316 3868
rect 259228 3816 259280 3868
rect 260656 3816 260708 3868
rect 261620 3816 261672 3868
rect 262956 3816 263008 3868
rect 263920 3816 263972 3868
rect 265348 3816 265400 3868
rect 268520 3816 268572 3868
rect 270040 3816 270092 3868
rect 270820 3816 270872 3868
rect 272432 3816 272484 3868
rect 275512 3816 275564 3868
rect 277124 3816 277176 3868
rect 277812 3816 277864 3868
rect 279516 3816 279568 3868
rect 284804 3816 284856 3868
rect 286600 3816 286652 3868
rect 292900 3816 292952 3868
rect 294880 3816 294932 3868
rect 299892 3816 299944 3868
rect 301964 3816 302016 3868
rect 306792 3816 306844 3868
rect 309048 3816 309100 3868
rect 572 3748 624 3800
rect 4112 3748 4164 3800
rect 7656 3748 7708 3800
rect 11012 3748 11064 3800
rect 12348 3748 12400 3800
rect 15704 3748 15756 3800
rect 15936 3748 15988 3800
rect 19108 3748 19160 3800
rect 21824 3748 21876 3800
rect 24904 3748 24956 3800
rect 25320 3748 25372 3800
rect 28400 3748 28452 3800
rect 31300 3748 31352 3800
rect 34196 3748 34248 3800
rect 34796 3748 34848 3800
rect 37692 3748 37744 3800
rect 40684 3748 40736 3800
rect 43488 3748 43540 3800
rect 44272 3748 44324 3800
rect 46984 3748 47036 3800
rect 47860 3748 47912 3800
rect 50480 3748 50532 3800
rect 51356 3748 51408 3800
rect 53976 3748 54028 3800
rect 54944 3748 54996 3800
rect 57380 3748 57432 3800
rect 58440 3748 58492 3800
rect 60876 3748 60928 3800
rect 64328 3748 64380 3800
rect 66672 3748 66724 3800
rect 67088 3748 67140 3800
rect 69064 3748 69116 3800
rect 70308 3748 70360 3800
rect 72468 3748 72520 3800
rect 73804 3748 73856 3800
rect 75964 3748 76016 3800
rect 79692 3748 79744 3800
rect 81760 3748 81812 3800
rect 86868 3748 86920 3800
rect 88752 3748 88804 3800
rect 95148 3748 95200 3800
rect 96848 3748 96900 3800
rect 103336 3748 103388 3800
rect 104944 3748 104996 3800
rect 216356 3748 216408 3800
rect 216864 3748 216916 3800
rect 222152 3748 222204 3800
rect 222752 3748 222804 3800
rect 224452 3748 224504 3800
rect 225144 3748 225196 3800
rect 230248 3748 230300 3800
rect 231032 3748 231084 3800
rect 231444 3748 231496 3800
rect 232228 3748 232280 3800
rect 232548 3748 232600 3800
rect 233424 3748 233476 3800
rect 233744 3748 233796 3800
rect 234620 3748 234672 3800
rect 237240 3748 237292 3800
rect 238116 3748 238168 3800
rect 238344 3748 238396 3800
rect 239312 3748 239364 3800
rect 239540 3748 239592 3800
rect 240508 3748 240560 3800
rect 240736 3748 240788 3800
rect 241704 3748 241756 3800
rect 241840 3748 241892 3800
rect 242900 3748 242952 3800
rect 245336 3748 245388 3800
rect 246396 3748 246448 3800
rect 246532 3748 246584 3800
rect 247592 3748 247644 3800
rect 250028 3748 250080 3800
rect 251180 3748 251232 3800
rect 252328 3748 252380 3800
rect 253480 3748 253532 3800
rect 255824 3748 255876 3800
rect 257068 3748 257120 3800
rect 258124 3748 258176 3800
rect 259460 3748 259512 3800
rect 260424 3748 260476 3800
rect 261760 3748 261812 3800
rect 262724 3748 262776 3800
rect 264152 3748 264204 3800
rect 265024 3748 265076 3800
rect 266544 3748 266596 3800
rect 267416 3748 267468 3800
rect 268844 3748 268896 3800
rect 269716 3748 269768 3800
rect 271236 3748 271288 3800
rect 272016 3748 272068 3800
rect 273628 3748 273680 3800
rect 276708 3748 276760 3800
rect 278320 3748 278372 3800
rect 279008 3748 279060 3800
rect 280712 3748 280764 3800
rect 283608 3748 283660 3800
rect 285404 3748 285456 3800
rect 287104 3748 287156 3800
rect 288992 3748 289044 3800
rect 291704 3748 291756 3800
rect 293684 3748 293736 3800
rect 294096 3748 294148 3800
rect 296076 3748 296128 3800
rect 298696 3748 298748 3800
rect 300768 3748 300820 3800
rect 300996 3748 301048 3800
rect 303160 3748 303212 3800
rect 307988 3748 308040 3800
rect 310244 3748 310296 3800
rect 316084 3748 316136 3800
rect 318524 3748 318576 3800
rect 323076 3748 323128 3800
rect 325608 3748 325660 3800
rect 6460 3000 6512 3052
rect 9864 3000 9916 3052
rect 63224 3000 63276 3052
rect 65524 3000 65576 3052
rect 535368 2932 535420 2984
rect 541992 2932 542044 2984
rect 573640 2932 573692 2984
rect 581000 2932 581052 2984
rect 18236 2864 18288 2916
rect 21456 2864 21508 2916
rect 253388 2864 253440 2916
rect 254676 2864 254728 2916
rect 506388 2864 506440 2916
rect 512460 2864 512512 2916
rect 516784 2864 516836 2916
rect 523040 2864 523092 2916
rect 524972 2864 525024 2916
rect 531320 2864 531372 2916
rect 536564 2864 536616 2916
rect 543188 2864 543240 2916
rect 544660 2864 544712 2916
rect 551468 2864 551520 2916
rect 553952 2864 554004 2916
rect 560852 2864 560904 2916
rect 574836 2864 574888 2916
rect 582196 2864 582248 2916
rect 4068 2796 4120 2848
rect 7472 2796 7524 2848
rect 9956 2796 10008 2848
rect 13268 2796 13320 2848
rect 17040 2796 17092 2848
rect 20260 2796 20312 2848
rect 28908 2796 28960 2848
rect 31852 2796 31904 2848
rect 35992 2796 36044 2848
rect 38844 2796 38896 2848
rect 39580 2796 39632 2848
rect 42340 2796 42392 2848
rect 62028 2796 62080 2848
rect 64420 2796 64472 2848
rect 65524 2796 65576 2848
rect 67824 2796 67876 2848
rect 248880 2796 248932 2848
rect 249984 2796 250036 2848
rect 251088 2796 251140 2848
rect 252376 2796 252428 2848
rect 254584 2796 254636 2848
rect 255872 2796 255924 2848
rect 309232 2796 309284 2848
rect 311440 2796 311492 2848
rect 315028 2796 315080 2848
rect 317328 2796 317380 2848
rect 411168 2796 411220 2848
rect 415492 2796 415544 2848
rect 440148 2796 440200 2848
rect 445024 2796 445076 2848
rect 449532 2796 449584 2848
rect 454500 2796 454552 2848
rect 478512 2796 478564 2848
rect 484032 2796 484084 2848
rect 487804 2796 487856 2848
rect 493508 2796 493560 2848
rect 507584 2796 507636 2848
rect 513564 2796 513616 2848
rect 515680 2796 515732 2848
rect 521844 2796 521896 2848
rect 545856 2796 545908 2848
rect 552664 2796 552716 2848
rect 3240 1300 3292 1352
rect 6368 1300 6420 1352
rect 60832 1300 60884 1352
rect 63316 1300 63368 1352
rect 67916 1300 67968 1352
rect 70124 1300 70176 1352
rect 76196 1300 76248 1352
rect 78220 1300 78272 1352
rect 83280 1300 83332 1352
rect 85212 1300 85264 1352
rect 85672 1300 85724 1352
rect 87512 1300 87564 1352
rect 89168 1300 89220 1352
rect 91008 1300 91060 1352
rect 91560 1300 91612 1352
rect 93308 1300 93360 1352
rect 93952 1300 94004 1352
rect 95700 1300 95752 1352
rect 97448 1300 97500 1352
rect 99104 1300 99156 1352
rect 101036 1300 101088 1352
rect 102600 1300 102652 1352
rect 104532 1300 104584 1352
rect 106096 1300 106148 1352
rect 106924 1300 106976 1352
rect 108396 1300 108448 1352
rect 109316 1300 109368 1352
rect 110696 1300 110748 1352
rect 112812 1300 112864 1352
rect 114192 1300 114244 1352
rect 116400 1300 116452 1352
rect 117688 1300 117740 1352
rect 119896 1300 119948 1352
rect 121184 1300 121236 1352
rect 125876 1300 125928 1352
rect 126980 1300 127032 1352
rect 129372 1300 129424 1352
rect 130476 1300 130528 1352
rect 130568 1300 130620 1352
rect 131580 1300 131632 1352
rect 131764 1300 131816 1352
rect 132776 1300 132828 1352
rect 132960 1300 133012 1352
rect 133972 1300 134024 1352
rect 137652 1300 137704 1352
rect 138572 1300 138624 1352
rect 144736 1300 144788 1352
rect 145564 1300 145616 1352
rect 145932 1300 145984 1352
rect 146668 1300 146720 1352
rect 148324 1300 148376 1352
rect 149060 1300 149112 1352
rect 154212 1300 154264 1352
rect 154856 1300 154908 1352
rect 162492 1300 162544 1352
rect 162952 1300 163004 1352
rect 266268 1300 266320 1352
rect 267740 1300 267792 1352
rect 273168 1300 273220 1352
rect 274824 1300 274876 1352
rect 280068 1300 280120 1352
rect 281908 1300 281960 1352
rect 282552 1300 282604 1352
rect 284300 1300 284352 1352
rect 288348 1300 288400 1352
rect 290188 1300 290240 1352
rect 295248 1300 295300 1352
rect 297272 1300 297324 1352
rect 297548 1300 297600 1352
rect 299664 1300 299716 1352
rect 302148 1300 302200 1352
rect 304356 1300 304408 1352
rect 305736 1300 305788 1352
rect 307944 1300 307996 1352
rect 310336 1300 310388 1352
rect 312636 1300 312688 1352
rect 313832 1300 313884 1352
rect 316224 1300 316276 1352
rect 317236 1300 317288 1352
rect 319720 1300 319772 1352
rect 321928 1300 321980 1352
rect 324412 1300 324464 1352
rect 325424 1300 325476 1352
rect 328000 1300 328052 1352
rect 328920 1300 328972 1352
rect 331588 1300 331640 1352
rect 332416 1300 332468 1352
rect 335084 1300 335136 1352
rect 335912 1300 335964 1352
rect 338672 1300 338724 1352
rect 339316 1300 339368 1352
rect 342168 1300 342220 1352
rect 345112 1300 345164 1352
rect 348056 1300 348108 1352
rect 349804 1300 349856 1352
rect 352840 1300 352892 1352
rect 353208 1300 353260 1352
rect 356336 1300 356388 1352
rect 356704 1300 356756 1352
rect 359924 1300 359976 1352
rect 362592 1300 362644 1352
rect 365812 1300 365864 1352
rect 367192 1300 367244 1352
rect 370596 1300 370648 1352
rect 370688 1300 370740 1352
rect 374092 1300 374144 1352
rect 376392 1300 376444 1352
rect 379980 1300 380032 1352
rect 385776 1300 385828 1352
rect 389456 1300 389508 1352
rect 395068 1300 395120 1352
rect 398932 1300 398984 1352
rect 399668 1300 399720 1352
rect 403624 1300 403676 1352
rect 405464 1300 405516 1352
rect 409604 1300 409656 1352
rect 413560 1300 413612 1352
rect 417884 1300 417936 1352
rect 422852 1300 422904 1352
rect 427268 1300 427320 1352
rect 427544 1300 427596 1352
rect 431868 1300 431920 1352
rect 433248 1300 433300 1352
rect 437848 1300 437900 1352
rect 442632 1300 442684 1352
rect 447416 1300 447468 1352
rect 448428 1300 448480 1352
rect 453304 1300 453356 1352
rect 458824 1300 458876 1352
rect 463976 1300 464028 1352
rect 468116 1300 468168 1352
rect 473084 1300 473136 1352
rect 475108 1300 475160 1352
rect 480536 1300 480588 1352
rect 485504 1300 485556 1352
rect 490748 1300 490800 1352
rect 497096 1300 497148 1352
rect 502984 1300 503036 1352
rect 504088 1300 504140 1352
rect 509700 1300 509752 1352
rect 513288 1300 513340 1352
rect 519544 1300 519596 1352
rect 526076 1300 526128 1352
rect 532148 1300 532200 1352
rect 534264 1300 534316 1352
rect 540428 1300 540480 1352
rect 541164 1300 541216 1352
rect 547880 1300 547932 1352
rect 548156 1300 548208 1352
rect 554780 1300 554832 1352
rect 555148 1300 555200 1352
rect 562048 1300 562100 1352
rect 566740 1300 566792 1352
rect 75000 1232 75052 1284
rect 77116 1232 77168 1284
rect 77392 1232 77444 1284
rect 79416 1232 79468 1284
rect 82084 1232 82136 1284
rect 84016 1232 84068 1284
rect 84476 1232 84528 1284
rect 86408 1232 86460 1284
rect 90364 1232 90416 1284
rect 92204 1232 92256 1284
rect 92756 1232 92808 1284
rect 94504 1232 94556 1284
rect 98644 1232 98696 1284
rect 100300 1232 100352 1284
rect 102232 1232 102284 1284
rect 103796 1232 103848 1284
rect 108120 1232 108172 1284
rect 109592 1232 109644 1284
rect 110512 1232 110564 1284
rect 111892 1232 111944 1284
rect 115204 1232 115256 1284
rect 116584 1232 116636 1284
rect 117596 1232 117648 1284
rect 118884 1232 118936 1284
rect 122288 1232 122340 1284
rect 123484 1232 123536 1284
rect 124680 1232 124732 1284
rect 125784 1232 125836 1284
rect 128176 1232 128228 1284
rect 129280 1232 129332 1284
rect 136456 1232 136508 1284
rect 137376 1232 137428 1284
rect 138848 1232 138900 1284
rect 139768 1232 139820 1284
rect 140044 1232 140096 1284
rect 140872 1232 140924 1284
rect 281356 1232 281408 1284
rect 283104 1232 283156 1284
rect 289452 1232 289504 1284
rect 291384 1232 291436 1284
rect 296444 1232 296496 1284
rect 298468 1232 298520 1284
rect 303344 1232 303396 1284
rect 305552 1232 305604 1284
rect 312544 1232 312596 1284
rect 315028 1232 315080 1284
rect 318432 1232 318484 1284
rect 320916 1232 320968 1284
rect 330024 1232 330076 1284
rect 332692 1232 332744 1284
rect 334716 1232 334768 1284
rect 337476 1232 337528 1284
rect 340512 1232 340564 1284
rect 343364 1232 343416 1284
rect 344008 1232 344060 1284
rect 346952 1232 347004 1284
rect 348608 1232 348660 1284
rect 351644 1232 351696 1284
rect 352104 1232 352156 1284
rect 355232 1232 355284 1284
rect 355600 1232 355652 1284
rect 358728 1232 358780 1284
rect 359096 1232 359148 1284
rect 362316 1232 362368 1284
rect 363696 1232 363748 1284
rect 367008 1232 367060 1284
rect 372988 1232 373040 1284
rect 376484 1232 376536 1284
rect 377588 1232 377640 1284
rect 381176 1232 381228 1284
rect 388076 1232 388128 1284
rect 391848 1232 391900 1284
rect 393872 1232 393924 1284
rect 397736 1232 397788 1284
rect 403164 1232 403216 1284
rect 407212 1232 407264 1284
rect 410064 1232 410116 1284
rect 414296 1232 414348 1284
rect 418252 1232 418304 1284
rect 422576 1232 422628 1284
rect 426348 1232 426400 1284
rect 430856 1232 430908 1284
rect 435640 1232 435692 1284
rect 439964 1232 440016 1284
rect 443736 1232 443788 1284
rect 448244 1232 448296 1284
rect 450728 1232 450780 1284
rect 455696 1232 455748 1284
rect 456524 1232 456576 1284
rect 461584 1232 461636 1284
rect 462228 1232 462280 1284
rect 467472 1232 467524 1284
rect 471612 1232 471664 1284
rect 476580 1232 476632 1284
rect 480904 1232 480956 1284
rect 486424 1232 486476 1284
rect 492496 1232 492548 1284
rect 498200 1232 498252 1284
rect 498292 1232 498344 1284
rect 503812 1232 503864 1284
rect 509884 1232 509936 1284
rect 515588 1232 515640 1284
rect 517980 1232 518032 1284
rect 523868 1232 523920 1284
rect 527272 1232 527324 1284
rect 533712 1232 533764 1284
rect 537668 1232 537720 1284
rect 544384 1232 544436 1284
rect 549352 1232 549404 1284
rect 556160 1232 556212 1284
rect 563244 1232 563296 1284
rect 570328 1232 570380 1284
rect 572536 1300 572588 1352
rect 579436 1300 579488 1352
rect 573548 1232 573600 1284
rect 576124 1232 576176 1284
rect 583392 1232 583444 1284
rect 99840 1164 99892 1216
rect 101496 1164 101548 1216
rect 114008 1164 114060 1216
rect 115388 1164 115440 1216
rect 311532 1164 311584 1216
rect 313832 1164 313884 1216
rect 319628 1164 319680 1216
rect 322112 1164 322164 1216
rect 327724 1164 327776 1216
rect 330392 1164 330444 1216
rect 331128 1164 331180 1216
rect 333888 1164 333940 1216
rect 337016 1164 337068 1216
rect 339868 1164 339920 1216
rect 341708 1164 341760 1216
rect 344560 1164 344612 1216
rect 357900 1164 357952 1216
rect 361120 1164 361172 1216
rect 364892 1164 364944 1216
rect 368204 1164 368256 1216
rect 375288 1164 375340 1216
rect 378876 1164 378928 1216
rect 381084 1164 381136 1216
rect 384764 1164 384816 1216
rect 390376 1164 390428 1216
rect 394240 1164 394292 1216
rect 396172 1164 396224 1216
rect 400128 1164 400180 1216
rect 400864 1164 400916 1216
rect 404820 1164 404872 1216
rect 407764 1164 407816 1216
rect 411904 1164 411956 1216
rect 420552 1164 420604 1216
rect 424968 1164 425020 1216
rect 425152 1164 425204 1216
rect 429660 1164 429712 1216
rect 441436 1164 441488 1216
rect 445852 1164 445904 1216
rect 447232 1164 447284 1216
rect 452108 1164 452160 1216
rect 454224 1164 454276 1216
rect 459192 1164 459244 1216
rect 460020 1164 460072 1216
rect 464804 1164 464856 1216
rect 470416 1164 470468 1216
rect 475752 1164 475804 1216
rect 477408 1164 477460 1216
rect 482468 1164 482520 1216
rect 483204 1164 483256 1216
rect 488816 1164 488868 1216
rect 490104 1164 490156 1216
rect 495532 1164 495584 1216
rect 505192 1164 505244 1216
rect 511264 1164 511316 1216
rect 514484 1164 514536 1216
rect 520372 1164 520424 1216
rect 521476 1164 521528 1216
rect 527824 1164 527876 1216
rect 528468 1164 528520 1216
rect 534540 1164 534592 1216
rect 542268 1164 542320 1216
rect 548708 1164 548760 1216
rect 556252 1164 556304 1216
rect 563152 1164 563204 1216
rect 569040 1164 569092 1216
rect 575940 1164 575992 1216
rect 5632 1096 5684 1148
rect 8668 1096 8720 1148
rect 111616 1096 111668 1148
rect 113088 1096 113140 1148
rect 123484 1096 123536 1148
rect 124772 1096 124824 1148
rect 320824 1096 320876 1148
rect 323308 1096 323360 1148
rect 360108 1096 360160 1148
rect 363512 1096 363564 1148
rect 382188 1096 382240 1148
rect 385960 1096 386012 1148
rect 389272 1096 389324 1148
rect 393044 1096 393096 1148
rect 398472 1096 398524 1148
rect 402520 1096 402572 1148
rect 404268 1096 404320 1148
rect 408408 1096 408460 1148
rect 408960 1096 409012 1148
rect 413100 1096 413152 1148
rect 415952 1096 416004 1148
rect 420184 1096 420236 1148
rect 429844 1096 429896 1148
rect 434444 1096 434496 1148
rect 436744 1096 436796 1148
rect 441528 1096 441580 1148
rect 446036 1096 446088 1148
rect 450912 1096 450964 1148
rect 457628 1096 457680 1148
rect 462412 1096 462464 1148
rect 464620 1096 464672 1148
rect 469864 1096 469916 1148
rect 472716 1096 472768 1148
rect 478144 1096 478196 1148
rect 486700 1096 486752 1148
rect 492312 1096 492364 1148
rect 500592 1096 500644 1148
rect 506480 1096 506532 1148
rect 510988 1096 511040 1148
rect 517152 1096 517204 1148
rect 522672 1096 522724 1148
rect 528652 1096 528704 1148
rect 530768 1096 530820 1148
rect 537208 1096 537260 1148
rect 543464 1096 543516 1148
rect 550272 1096 550324 1148
rect 550456 1096 550508 1148
rect 556988 1096 557040 1148
rect 558552 1096 558604 1148
rect 565268 1096 565320 1148
rect 567844 1096 567896 1148
rect 575112 1096 575164 1148
rect 378784 1028 378836 1080
rect 382372 1028 382424 1080
rect 386880 1028 386932 1080
rect 390652 1028 390704 1080
rect 417056 1028 417108 1080
rect 421380 1028 421432 1080
rect 428648 1028 428700 1080
rect 433248 1028 433300 1080
rect 437940 1028 437992 1080
rect 442632 1028 442684 1080
rect 455328 1028 455380 1080
rect 460020 1028 460072 1080
rect 465816 1028 465868 1080
rect 470692 1028 470744 1080
rect 473912 1028 473964 1080
rect 478972 1028 479024 1080
rect 482008 1028 482060 1080
rect 487252 1028 487304 1080
rect 491208 1028 491260 1080
rect 497096 1028 497148 1080
rect 499396 1028 499448 1080
rect 505376 1028 505428 1080
rect 508688 1028 508740 1080
rect 514760 1028 514812 1080
rect 519176 1028 519228 1080
rect 525432 1028 525484 1080
rect 531872 1028 531924 1080
rect 538220 1028 538272 1080
rect 538864 1028 538916 1080
rect 545488 1028 545540 1080
rect 546960 1028 547012 1080
rect 553768 1028 553820 1080
rect 560944 1028 560996 1080
rect 567660 1028 567712 1080
rect 571248 1028 571300 1080
rect 578608 1028 578660 1080
rect 326620 960 326672 1012
rect 329196 960 329248 1012
rect 374184 960 374236 1012
rect 377680 960 377732 1012
rect 379888 960 379940 1012
rect 383568 960 383620 1012
rect 414756 960 414808 1012
rect 418988 960 419040 1012
rect 424048 960 424100 1012
rect 428464 960 428516 1012
rect 432144 960 432196 1012
rect 436744 960 436796 1012
rect 439136 960 439188 1012
rect 443828 960 443880 1012
rect 453028 960 453080 1012
rect 458088 960 458140 1012
rect 466920 960 466972 1012
rect 472256 960 472308 1012
rect 476212 960 476264 1012
rect 481364 960 481416 1012
rect 489000 960 489052 1012
rect 494704 960 494756 1012
rect 494796 960 494848 1012
rect 500592 960 500644 1012
rect 501788 960 501840 1012
rect 507308 960 507360 1012
rect 512184 960 512236 1012
rect 517980 960 518032 1012
rect 523776 960 523828 1012
rect 529940 960 529992 1012
rect 533068 960 533120 1012
rect 539600 960 539652 1012
rect 540060 960 540112 1012
rect 546500 960 546552 1012
rect 551652 960 551704 1012
rect 558552 960 558604 1012
rect 561956 960 562008 1012
rect 568764 960 568816 1012
rect 570144 960 570196 1012
rect 577044 960 577096 1012
rect 8760 892 8812 944
rect 12164 892 12216 944
rect 121092 892 121144 944
rect 122380 892 122432 944
rect 463424 892 463476 944
rect 468300 892 468352 944
rect 479708 892 479760 944
rect 484860 892 484912 944
rect 493600 892 493652 944
rect 499396 892 499448 944
rect 502892 892 502944 944
rect 508872 892 508924 944
rect 520188 892 520240 944
rect 526260 892 526312 944
rect 529572 892 529624 944
rect 536104 892 536156 944
rect 559656 892 559708 944
rect 566832 892 566884 944
rect 347504 824 347556 876
rect 350448 824 350500 876
rect 361396 824 361448 876
rect 364616 824 364668 876
rect 368388 824 368440 876
rect 371700 824 371752 876
rect 371792 824 371844 876
rect 375288 824 375340 876
rect 384580 824 384632 876
rect 388260 824 388312 876
rect 391572 824 391624 876
rect 395344 824 395396 876
rect 397368 824 397420 876
rect 401324 824 401376 876
rect 406660 824 406712 876
rect 410800 824 410852 876
rect 419356 824 419408 876
rect 423404 824 423456 876
rect 434352 824 434404 876
rect 439136 824 439188 876
rect 444932 824 444984 876
rect 449808 824 449860 876
rect 461124 824 461176 876
rect 466276 824 466328 876
rect 484308 824 484360 876
rect 489920 824 489972 876
rect 495992 824 496044 876
rect 501788 824 501840 876
rect 552756 824 552808 876
rect 559748 824 559800 876
rect 52552 688 52604 740
rect 55036 688 55088 740
rect 59636 688 59688 740
rect 61936 688 61988 740
rect 105728 688 105780 740
rect 107292 688 107344 740
rect 274364 688 274416 740
rect 276020 688 276072 740
rect 333520 688 333572 740
rect 336280 688 336332 740
rect 338212 688 338264 740
rect 340972 688 341024 740
rect 342812 688 342864 740
rect 345756 688 345808 740
rect 346308 688 346360 740
rect 349252 688 349304 740
rect 350908 688 350960 740
rect 354036 688 354088 740
rect 365996 688 366048 740
rect 369400 688 369452 740
rect 369492 688 369544 740
rect 372896 688 372948 740
rect 451832 688 451884 740
rect 456524 688 456576 740
rect 69112 552 69164 604
rect 71320 552 71372 604
rect 290648 552 290700 604
rect 292580 552 292632 604
rect 304540 552 304592 604
rect 306748 552 306800 604
rect 324228 552 324280 604
rect 326804 552 326856 604
rect 416688 552 416740 604
rect 557540 552 557592 604
rect 564440 552 564492 604
rect 412456 348 412508 400
rect 565452 416 565504 468
rect 572904 416 572956 468
rect 401968 144 402020 196
rect 406200 144 406252 196
rect 383384 76 383436 128
rect 386788 76 386840 128
rect 421748 76 421800 128
rect 425796 76 425848 128
rect 354404 8 354456 60
rect 357348 8 357400 60
rect 392676 8 392728 60
rect 396172 8 396224 60
rect 431040 8 431092 60
rect 435180 8 435232 60
rect 469312 8 469364 60
rect 474188 8 474240 60
rect 564256 8 564308 60
rect 571340 8 571392 60
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700806 8156 703520
rect 3884 700800 3936 700806
rect 3884 700742 3936 700748
rect 8116 700800 8168 700806
rect 8116 700742 8168 700748
rect 18 698184 74 698193
rect 18 698119 74 698128
rect 32 684593 60 698119
rect 3896 697966 3924 700742
rect 24320 700262 24348 703520
rect 40512 700262 40540 703520
rect 72988 700262 73016 703520
rect 89180 700262 89208 703520
rect 105464 700330 105492 703520
rect 105452 700324 105504 700330
rect 105452 700266 105504 700272
rect 113916 700324 113968 700330
rect 113916 700266 113968 700272
rect 24308 700256 24360 700262
rect 24308 700198 24360 700204
rect 25964 700256 26016 700262
rect 25964 700198 26016 700204
rect 40500 700256 40552 700262
rect 40500 700198 40552 700204
rect 47952 700256 48004 700262
rect 47952 700198 48004 700204
rect 70032 700256 70084 700262
rect 70032 700198 70084 700204
rect 72976 700256 73028 700262
rect 72976 700198 73028 700204
rect 89168 700256 89220 700262
rect 89168 700198 89220 700204
rect 91928 700256 91980 700262
rect 91928 700198 91980 700204
rect 25976 698170 26004 700198
rect 47964 698170 47992 700198
rect 70044 698170 70072 700198
rect 25976 698142 26048 698170
rect 47964 698142 48036 698170
rect 3896 697938 4046 697966
rect 26020 697959 26048 698142
rect 48008 697959 48036 698142
rect 69996 698142 70072 698170
rect 91940 698170 91968 700198
rect 113928 698170 113956 700266
rect 137848 700262 137876 703520
rect 154132 700262 154160 703520
rect 170324 700330 170352 703520
rect 170312 700324 170364 700330
rect 170312 700266 170364 700272
rect 179880 700324 179932 700330
rect 179880 700266 179932 700272
rect 135996 700256 136048 700262
rect 135996 700198 136048 700204
rect 137836 700256 137888 700262
rect 137836 700198 137888 700204
rect 154120 700256 154172 700262
rect 154120 700198 154172 700204
rect 157892 700256 157944 700262
rect 157892 700198 157944 700204
rect 136008 698170 136036 700198
rect 91940 698142 92012 698170
rect 113928 698142 114000 698170
rect 69996 697959 70024 698142
rect 91984 697959 92012 698142
rect 113972 697959 114000 698142
rect 135960 698142 136036 698170
rect 157904 698170 157932 700198
rect 179892 698170 179920 700266
rect 202800 700262 202828 703520
rect 218992 700330 219020 703520
rect 235184 700330 235212 703520
rect 218980 700324 219032 700330
rect 218980 700266 219032 700272
rect 223856 700324 223908 700330
rect 223856 700266 223908 700272
rect 235172 700324 235224 700330
rect 235172 700266 235224 700272
rect 245844 700324 245896 700330
rect 245844 700266 245896 700272
rect 201960 700256 202012 700262
rect 201960 700198 202012 700204
rect 202788 700256 202840 700262
rect 202788 700198 202840 700204
rect 201972 698170 202000 700198
rect 157904 698142 157976 698170
rect 179892 698142 179964 698170
rect 135960 697959 135988 698142
rect 157948 697959 157976 698142
rect 179936 697959 179964 698142
rect 201924 698142 202000 698170
rect 223868 698170 223896 700266
rect 245856 698170 245884 700266
rect 267660 699802 267688 703520
rect 283852 700330 283880 703520
rect 300136 700330 300164 703520
rect 283840 700324 283892 700330
rect 283840 700266 283892 700272
rect 289820 700324 289872 700330
rect 289820 700266 289872 700272
rect 300124 700324 300176 700330
rect 300124 700266 300176 700272
rect 311900 700324 311952 700330
rect 311900 700266 311952 700272
rect 267660 699774 267872 699802
rect 267844 698170 267872 699774
rect 289832 698170 289860 700266
rect 311912 698170 311940 700266
rect 332520 700126 332548 703520
rect 348804 700602 348832 703520
rect 348792 700596 348844 700602
rect 348792 700538 348844 700544
rect 355876 700596 355928 700602
rect 355876 700538 355928 700544
rect 332508 700120 332560 700126
rect 332508 700062 332560 700068
rect 333888 700120 333940 700126
rect 333888 700062 333940 700068
rect 333900 698170 333928 700062
rect 355888 698170 355916 700538
rect 364996 700330 365024 703520
rect 364984 700324 365036 700330
rect 364984 700266 365036 700272
rect 377864 700324 377916 700330
rect 377864 700266 377916 700272
rect 377876 698170 377904 700266
rect 397472 700262 397500 703520
rect 413664 700262 413692 703520
rect 429856 700330 429884 703520
rect 429844 700324 429896 700330
rect 429844 700266 429896 700272
rect 443828 700324 443880 700330
rect 443828 700266 443880 700272
rect 397460 700256 397512 700262
rect 397460 700198 397512 700204
rect 399852 700256 399904 700262
rect 399852 700198 399904 700204
rect 413652 700256 413704 700262
rect 413652 700198 413704 700204
rect 421840 700256 421892 700262
rect 421840 700198 421892 700204
rect 399864 698170 399892 700198
rect 421852 698170 421880 700198
rect 443840 698170 443868 700266
rect 462332 700262 462360 703520
rect 478524 700330 478552 703520
rect 494808 700330 494836 703520
rect 527192 700330 527220 703520
rect 543476 700330 543504 703520
rect 559668 700330 559696 703520
rect 478512 700324 478564 700330
rect 478512 700266 478564 700272
rect 487804 700324 487856 700330
rect 487804 700266 487856 700272
rect 494796 700324 494848 700330
rect 494796 700266 494848 700272
rect 509792 700324 509844 700330
rect 509792 700266 509844 700272
rect 527180 700324 527232 700330
rect 527180 700266 527232 700272
rect 531780 700324 531832 700330
rect 531780 700266 531832 700272
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 553768 700324 553820 700330
rect 553768 700266 553820 700272
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 575756 700324 575808 700330
rect 575756 700266 575808 700272
rect 462320 700256 462372 700262
rect 462320 700198 462372 700204
rect 465816 700256 465868 700262
rect 465816 700198 465868 700204
rect 465828 698170 465856 700198
rect 487816 698170 487844 700266
rect 509804 698170 509832 700266
rect 531792 698170 531820 700266
rect 553780 698170 553808 700266
rect 575768 698170 575796 700266
rect 223868 698142 223940 698170
rect 245856 698142 245928 698170
rect 267844 698142 267916 698170
rect 289832 698142 289904 698170
rect 311912 698142 311984 698170
rect 333900 698142 333972 698170
rect 355888 698142 355960 698170
rect 377876 698142 377948 698170
rect 399864 698142 399936 698170
rect 421852 698142 421924 698170
rect 443840 698142 443912 698170
rect 465828 698142 465900 698170
rect 487816 698142 487888 698170
rect 509804 698142 509876 698170
rect 531792 698142 531864 698170
rect 553780 698142 553852 698170
rect 575768 698142 575840 698170
rect 201924 697959 201952 698142
rect 223912 697959 223940 698142
rect 245900 697959 245928 698142
rect 267888 697959 267916 698142
rect 289876 697959 289904 698142
rect 311956 697959 311984 698142
rect 333944 697959 333972 698142
rect 355932 697959 355960 698142
rect 377920 697959 377948 698142
rect 399908 697959 399936 698142
rect 421896 697959 421924 698142
rect 443884 697959 443912 698142
rect 465872 697959 465900 698142
rect 487860 697959 487888 698142
rect 509848 697959 509876 698142
rect 531836 697959 531864 698142
rect 553824 697959 553852 698142
rect 575812 697959 575840 698142
rect 18 684584 74 684593
rect 18 684519 74 684528
rect 579986 683904 580042 683913
rect 579986 683839 580042 683848
rect 580000 682514 580028 683839
rect 578424 682508 578476 682514
rect 578424 682450 578476 682456
rect 579988 682508 580040 682514
rect 579988 682450 580040 682456
rect 578436 682281 578464 682450
rect 578422 682272 578478 682281
rect 578422 682207 578478 682216
rect 2778 681048 2834 681057
rect 2778 680983 2834 680992
rect 2792 671265 2820 680983
rect 2778 671256 2834 671265
rect 2778 671191 2834 671200
rect 579526 670712 579582 670721
rect 579526 670647 579582 670656
rect 579540 666505 579568 670647
rect 579526 666496 579582 666505
rect 579526 666431 579582 666440
rect 3422 664060 3478 664069
rect 3422 663995 3478 664004
rect 3436 658209 3464 663995
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 578882 650720 578938 650729
rect 578882 650655 578938 650664
rect 18 647048 74 647057
rect 18 646983 74 646992
rect 32 632641 60 646983
rect 578896 644065 578924 650655
rect 578882 644056 578938 644065
rect 578882 643991 578938 644000
rect 579526 634944 579582 634953
rect 579526 634879 579582 634888
rect 579540 634814 579568 634879
rect 579540 634786 579660 634814
rect 18 632632 74 632641
rect 18 632567 74 632576
rect 579632 630873 579660 634786
rect 579618 630864 579674 630873
rect 579618 630799 579674 630808
rect 2778 630320 2834 630329
rect 2778 630255 2834 630264
rect 2792 619177 2820 630255
rect 2778 619168 2834 619177
rect 2778 619103 2834 619112
rect 579526 619168 579582 619177
rect 579582 619126 579660 619154
rect 579526 619103 579582 619112
rect 579632 617545 579660 619126
rect 579618 617536 579674 617545
rect 579618 617471 579674 617480
rect 3422 613308 3478 613317
rect 3422 613243 3478 613252
rect 3436 606121 3464 613243
rect 3422 606112 3478 606121
rect 3422 606047 3478 606056
rect 578882 603392 578938 603401
rect 578882 603327 578938 603336
rect 18 596320 74 596329
rect 18 596255 74 596264
rect 32 580553 60 596255
rect 578896 591025 578924 603327
rect 578882 591016 578938 591025
rect 578882 590951 578938 590960
rect 578882 587616 578938 587625
rect 578882 587551 578938 587560
rect 18 580544 74 580553
rect 18 580479 74 580488
rect 18 579456 74 579465
rect 18 579391 74 579400
rect 32 567225 60 579391
rect 578896 577697 578924 587551
rect 578882 577688 578938 577697
rect 578882 577623 578938 577632
rect 578882 571840 578938 571849
rect 578882 571775 578938 571784
rect 18 567216 74 567225
rect 18 567151 74 567160
rect 578896 564369 578924 571775
rect 578882 564360 578938 564369
rect 578882 564295 578938 564304
rect 2778 562592 2834 562601
rect 2778 562527 2834 562536
rect 2792 553897 2820 562527
rect 578882 556064 578938 556073
rect 578882 555999 578938 556008
rect 2778 553888 2834 553897
rect 2778 553823 2834 553832
rect 18 545592 74 545601
rect 18 545527 74 545536
rect 32 528193 60 545527
rect 578896 537849 578924 555999
rect 578974 540288 579030 540297
rect 578974 540223 579030 540232
rect 578882 537840 578938 537849
rect 578882 537775 578938 537784
rect 110 528592 166 528601
rect 110 528527 166 528536
rect 18 528184 74 528193
rect 18 528119 74 528128
rect 124 515409 152 528527
rect 578882 524648 578938 524657
rect 578882 524583 578938 524592
rect 110 515400 166 515409
rect 110 515335 166 515344
rect 2778 511864 2834 511873
rect 2778 511799 2834 511808
rect 2792 501809 2820 511799
rect 578896 511329 578924 524583
rect 578988 524521 579016 540223
rect 578974 524512 579030 524521
rect 578974 524447 579030 524456
rect 578882 511320 578938 511329
rect 578882 511255 578938 511264
rect 578882 508736 578938 508745
rect 578882 508671 578938 508680
rect 2778 501800 2834 501809
rect 2778 501735 2834 501744
rect 18 494864 74 494873
rect 18 494799 74 494808
rect 32 476105 60 494799
rect 578896 484673 578924 508671
rect 578974 492824 579030 492833
rect 578974 492759 579030 492768
rect 578882 484664 578938 484673
rect 578882 484599 578938 484608
rect 110 477864 166 477873
rect 110 477799 166 477808
rect 18 476096 74 476105
rect 18 476031 74 476040
rect 124 463185 152 477799
rect 578988 471481 579016 492759
rect 579066 477320 579122 477329
rect 579066 477255 579122 477264
rect 578974 471472 579030 471481
rect 578974 471407 579030 471416
rect 110 463176 166 463185
rect 110 463111 166 463120
rect 578882 461544 578938 461553
rect 578882 461479 578938 461488
rect 18 461000 74 461009
rect 18 460935 74 460944
rect 32 449857 60 460935
rect 18 449848 74 449857
rect 18 449783 74 449792
rect 18 444136 74 444145
rect 18 444071 74 444080
rect 32 423638 60 444071
rect 578896 431633 578924 461479
rect 579080 458153 579108 477255
rect 579066 458144 579122 458153
rect 579066 458079 579122 458088
rect 578974 445632 579030 445641
rect 578974 445567 579030 445576
rect 578882 431624 578938 431633
rect 578882 431559 578938 431568
rect 110 427136 166 427145
rect 110 427071 166 427080
rect 20 423632 72 423638
rect 20 423574 72 423580
rect 124 411097 152 427071
rect 572 423632 624 423638
rect 570 423600 572 423609
rect 624 423600 626 423609
rect 570 423535 626 423544
rect 578988 418305 579016 445567
rect 579066 429856 579122 429865
rect 579066 429791 579122 429800
rect 578974 418296 579030 418305
rect 578974 418231 579030 418240
rect 578882 414216 578938 414225
rect 578882 414151 578938 414160
rect 110 411088 166 411097
rect 110 411023 166 411032
rect 294 410136 350 410145
rect 294 410071 350 410080
rect 308 398041 336 410071
rect 578238 398440 578294 398449
rect 578238 398375 578294 398384
rect 294 398032 350 398041
rect 294 397967 350 397976
rect 578252 397526 578280 398375
rect 578240 397520 578292 397526
rect 578240 397462 578292 397468
rect 18 393408 74 393417
rect 18 393343 74 393352
rect 32 371929 60 393343
rect 578896 378457 578924 414151
rect 579080 404977 579108 429791
rect 579066 404968 579122 404977
rect 579066 404903 579122 404912
rect 580264 397520 580316 397526
rect 580264 397462 580316 397468
rect 578974 382528 579030 382537
rect 578974 382463 579030 382472
rect 578882 378448 578938 378457
rect 578882 378383 578938 378392
rect 110 376408 166 376417
rect 110 376343 166 376352
rect 18 371920 74 371929
rect 18 371855 74 371864
rect 18 359408 74 359417
rect 18 359343 74 359352
rect 32 345953 60 359343
rect 124 358737 152 376343
rect 578882 366888 578938 366897
rect 578882 366823 578938 366832
rect 110 358728 166 358737
rect 110 358663 166 358672
rect 578330 351112 578386 351121
rect 578330 351047 578332 351056
rect 578384 351047 578386 351056
rect 578332 351018 578384 351024
rect 18 345944 74 345953
rect 18 345879 74 345888
rect 18 342544 74 342553
rect 18 342479 74 342488
rect 32 319841 60 342479
rect 110 325680 166 325689
rect 110 325615 166 325624
rect 18 319832 74 319841
rect 18 319767 74 319776
rect 18 308680 74 308689
rect 18 308615 74 308624
rect 32 293729 60 308615
rect 124 306513 152 325615
rect 578896 325281 578924 366823
rect 578988 351937 579016 382463
rect 580276 365129 580304 397462
rect 580262 365120 580318 365129
rect 580262 365055 580318 365064
rect 578974 351928 579030 351937
rect 578974 351863 579030 351872
rect 580264 351076 580316 351082
rect 580264 351018 580316 351024
rect 578974 335472 579030 335481
rect 578974 335407 579030 335416
rect 578882 325272 578938 325281
rect 578882 325207 578938 325216
rect 578882 319560 578938 319569
rect 578882 319495 578938 319504
rect 110 306504 166 306513
rect 110 306439 166 306448
rect 578514 303784 578570 303793
rect 578514 303719 578516 303728
rect 578568 303719 578570 303728
rect 578516 303690 578568 303696
rect 18 293720 74 293729
rect 18 293655 74 293664
rect 18 291816 74 291825
rect 18 291751 74 291760
rect 32 267481 60 291751
rect 110 274816 166 274825
rect 110 274751 166 274760
rect 18 267472 74 267481
rect 18 267407 74 267416
rect 124 254697 152 274751
rect 578896 273222 578924 319495
rect 578988 298761 579016 335407
rect 580276 312089 580304 351018
rect 580262 312080 580318 312089
rect 580262 312015 580318 312024
rect 580264 303748 580316 303754
rect 580264 303690 580316 303696
rect 578974 298752 579030 298761
rect 578974 298687 579030 298696
rect 578974 288008 579030 288017
rect 578974 287943 579030 287952
rect 578884 273216 578936 273222
rect 578884 273158 578936 273164
rect 202 257952 258 257961
rect 202 257887 258 257896
rect 110 254688 166 254697
rect 110 254623 166 254632
rect 216 241505 244 257887
rect 578606 256456 578662 256465
rect 578606 256391 578662 256400
rect 578620 255338 578648 256391
rect 578608 255332 578660 255338
rect 578608 255274 578660 255280
rect 578988 245585 579016 287943
rect 579066 272232 579122 272241
rect 579066 272167 579122 272176
rect 578974 245576 579030 245585
rect 578974 245511 579030 245520
rect 202 241496 258 241505
rect 202 241431 258 241440
rect 18 240816 74 240825
rect 18 240751 74 240760
rect 32 215257 60 240751
rect 578882 240680 578938 240689
rect 578882 240615 578938 240624
rect 110 224088 166 224097
rect 110 224023 166 224032
rect 18 215248 74 215257
rect 18 215183 74 215192
rect 124 202473 152 224023
rect 578330 209264 578386 209273
rect 578330 209199 578386 209208
rect 578344 208418 578372 209199
rect 578332 208412 578384 208418
rect 578332 208354 578384 208360
rect 202 207224 258 207233
rect 202 207159 258 207168
rect 110 202464 166 202473
rect 110 202399 166 202408
rect 18 190224 74 190233
rect 18 190159 74 190168
rect 32 163441 60 190159
rect 216 189145 244 207159
rect 578896 205737 578924 240615
rect 579080 232393 579108 272167
rect 580276 258913 580304 303690
rect 580816 273216 580868 273222
rect 580816 273158 580868 273164
rect 580828 272241 580856 273158
rect 580814 272232 580870 272241
rect 580814 272167 580870 272176
rect 580262 258904 580318 258913
rect 580262 258839 580318 258848
rect 580264 255332 580316 255338
rect 580264 255274 580316 255280
rect 579066 232384 579122 232393
rect 579066 232319 579122 232328
rect 578974 225040 579030 225049
rect 578974 224975 579030 224984
rect 578882 205728 578938 205737
rect 578882 205663 578938 205672
rect 578882 193352 578938 193361
rect 578882 193287 578938 193296
rect 202 189136 258 189145
rect 202 189071 258 189080
rect 110 173360 166 173369
rect 110 173295 166 173304
rect 18 163432 74 163441
rect 18 163367 74 163376
rect 124 150385 152 173295
rect 578896 165889 578924 193287
rect 578988 192545 579016 224975
rect 580276 219065 580304 255274
rect 580262 219056 580318 219065
rect 580262 218991 580318 219000
rect 580264 208412 580316 208418
rect 580264 208354 580316 208360
rect 578974 192536 579030 192545
rect 578974 192471 579030 192480
rect 580276 179217 580304 208354
rect 580262 179208 580318 179217
rect 580262 179143 580318 179152
rect 578974 177576 579030 177585
rect 578974 177511 579030 177520
rect 578882 165880 578938 165889
rect 578882 165815 578938 165824
rect 578882 161936 578938 161945
rect 578882 161871 578938 161880
rect 202 156360 258 156369
rect 202 156295 258 156304
rect 110 150376 166 150385
rect 110 150311 166 150320
rect 18 139496 74 139505
rect 18 139431 74 139440
rect 32 111217 60 139431
rect 216 137329 244 156295
rect 578896 139369 578924 161871
rect 578988 152697 579016 177511
rect 578974 152688 579030 152697
rect 578974 152623 579030 152632
rect 578974 146160 579030 146169
rect 578974 146095 579030 146104
rect 578882 139360 578938 139369
rect 578882 139295 578938 139304
rect 202 137320 258 137329
rect 202 137255 258 137264
rect 578882 130248 578938 130257
rect 578882 130183 578938 130192
rect 110 122496 166 122505
rect 110 122431 166 122440
rect 18 111208 74 111217
rect 18 111143 74 111152
rect 18 105632 74 105641
rect 18 105567 74 105576
rect 32 85241 60 105567
rect 124 97889 152 122431
rect 578896 112849 578924 130183
rect 578988 126041 579016 146095
rect 578974 126032 579030 126041
rect 578974 125967 579030 125976
rect 578974 114608 579030 114617
rect 578974 114543 579030 114552
rect 578882 112840 578938 112849
rect 578882 112775 578938 112784
rect 578988 99521 579016 114543
rect 578974 99512 579030 99521
rect 578974 99447 579030 99456
rect 578882 98832 578938 98841
rect 578882 98767 578938 98776
rect 110 97880 166 97889
rect 110 97815 166 97824
rect 110 88768 166 88777
rect 110 88703 166 88712
rect 18 85232 74 85241
rect 18 85167 74 85176
rect 124 71913 152 88703
rect 578896 86193 578924 98767
rect 578882 86184 578938 86193
rect 578882 86119 578938 86128
rect 578882 83056 578938 83065
rect 578882 82991 578938 83000
rect 578896 73001 578924 82991
rect 578882 72992 578938 73001
rect 578882 72927 578938 72936
rect 110 71904 166 71913
rect 110 71839 166 71848
rect 294 71360 350 71369
rect 294 71295 350 71304
rect 308 59129 336 71295
rect 578238 67280 578294 67289
rect 578238 67215 578294 67224
rect 578252 60722 578280 67215
rect 578240 60716 578292 60722
rect 578240 60658 578292 60664
rect 580816 60716 580868 60722
rect 580816 60658 580868 60664
rect 580828 59673 580856 60658
rect 580814 59664 580870 59673
rect 580814 59599 580870 59608
rect 294 59120 350 59129
rect 294 59055 350 59064
rect 2778 54904 2834 54913
rect 2778 54839 2834 54848
rect 2792 45529 2820 54839
rect 579526 51504 579582 51513
rect 579526 51439 579582 51448
rect 579540 46345 579568 51439
rect 579526 46336 579582 46345
rect 579526 46271 579582 46280
rect 2778 45520 2834 45529
rect 2778 45455 2834 45464
rect 2042 37904 2098 37913
rect 2042 37839 2098 37848
rect 2056 32473 2084 37839
rect 579526 35728 579582 35737
rect 579582 35686 579660 35714
rect 579526 35663 579582 35672
rect 579632 33153 579660 35686
rect 579618 33144 579674 33153
rect 579618 33079 579674 33088
rect 2042 32464 2098 32473
rect 2042 32399 2098 32408
rect 1306 21040 1362 21049
rect 1306 20975 1362 20984
rect 1320 19417 1348 20975
rect 1306 19408 1362 19417
rect 1306 19343 1362 19352
rect 579618 6624 579674 6633
rect 579618 6559 579674 6568
rect 2778 6488 2834 6497
rect 2778 6423 2834 6432
rect 2792 4185 2820 6423
rect 2778 4176 2834 4185
rect 2778 4111 2834 4120
rect 579526 4176 579582 4185
rect 579632 4162 579660 6559
rect 579582 4134 579660 4162
rect 579526 4111 579582 4120
rect 1676 3868 1728 3874
rect 1676 3810 1728 3816
rect 572 3800 624 3806
rect 572 3742 624 3748
rect 584 480 612 3742
rect 1688 480 1716 3810
rect 4124 3806 4152 4012
rect 5228 3874 5256 4012
rect 5216 3868 5268 3874
rect 5216 3810 5268 3816
rect 4112 3800 4164 3806
rect 6424 3754 6452 4012
rect 7528 3754 7556 4012
rect 4112 3742 4164 3748
rect 6380 3726 6452 3754
rect 7484 3726 7556 3754
rect 7656 3800 7708 3806
rect 8724 3754 8752 4012
rect 9920 3754 9948 4012
rect 11024 3806 11052 4012
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 7656 3742 7708 3748
rect 4068 2848 4120 2854
rect 4068 2790 4120 2796
rect 3240 1352 3292 1358
rect 3240 1294 3292 1300
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 354 2954 480
rect 3252 354 3280 1294
rect 4080 480 4108 2790
rect 6380 1358 6408 3726
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 6368 1352 6420 1358
rect 6368 1294 6420 1300
rect 5632 1148 5684 1154
rect 5632 1090 5684 1096
rect 2842 326 3280 354
rect 2842 -960 2954 326
rect 4038 -960 4150 480
rect 5234 354 5346 480
rect 5644 354 5672 1090
rect 6472 480 6500 2994
rect 7484 2854 7512 3726
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 7668 480 7696 3742
rect 8680 3726 8752 3754
rect 9876 3726 9948 3754
rect 11012 3800 11064 3806
rect 11012 3742 11064 3748
rect 8680 1154 8708 3726
rect 9876 3058 9904 3726
rect 9864 3052 9916 3058
rect 9864 2994 9916 3000
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 8668 1148 8720 1154
rect 8668 1090 8720 1096
rect 8760 944 8812 950
rect 8760 886 8812 892
rect 8772 480 8800 886
rect 9968 480 9996 2790
rect 11164 480 11192 3878
rect 12220 3754 12248 4012
rect 12176 3726 12248 3754
rect 12348 3800 12400 3806
rect 13324 3754 13352 4012
rect 14520 3942 14548 4012
rect 14508 3936 14560 3942
rect 14508 3878 14560 3884
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 13544 3868 13596 3874
rect 13544 3810 13596 3816
rect 12348 3742 12400 3748
rect 12176 950 12204 3726
rect 12164 944 12216 950
rect 12164 886 12216 892
rect 12360 480 12388 3742
rect 13280 3726 13352 3754
rect 13280 2854 13308 3726
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 13556 480 13584 3810
rect 14752 480 14780 3878
rect 15716 3806 15744 4012
rect 16820 3874 16848 4012
rect 18016 3942 18044 4012
rect 18004 3936 18056 3942
rect 18004 3878 18056 3884
rect 16808 3868 16860 3874
rect 16808 3810 16860 3816
rect 19120 3806 19148 4012
rect 19432 3868 19484 3874
rect 19432 3810 19484 3816
rect 15704 3800 15756 3806
rect 15704 3742 15756 3748
rect 15936 3800 15988 3806
rect 15936 3742 15988 3748
rect 19108 3800 19160 3806
rect 19108 3742 19160 3748
rect 15948 480 15976 3742
rect 18236 2916 18288 2922
rect 18236 2858 18288 2864
rect 17040 2848 17092 2854
rect 17040 2790 17092 2796
rect 17052 480 17080 2790
rect 18248 480 18276 2858
rect 19444 480 19472 3810
rect 20316 3754 20344 4012
rect 20628 3936 20680 3942
rect 20628 3878 20680 3884
rect 20272 3726 20344 3754
rect 20272 2854 20300 3726
rect 20260 2848 20312 2854
rect 20260 2790 20312 2796
rect 20640 480 20668 3878
rect 21512 3754 21540 4012
rect 22616 3874 22644 4012
rect 23812 3942 23840 4012
rect 23800 3936 23852 3942
rect 23800 3878 23852 3884
rect 24216 3936 24268 3942
rect 24216 3878 24268 3884
rect 22604 3868 22656 3874
rect 22604 3810 22656 3816
rect 23020 3868 23072 3874
rect 23020 3810 23072 3816
rect 21468 3726 21540 3754
rect 21824 3800 21876 3806
rect 21824 3742 21876 3748
rect 21468 2922 21496 3726
rect 21456 2916 21508 2922
rect 21456 2858 21508 2864
rect 21836 480 21864 3742
rect 23032 480 23060 3810
rect 24228 480 24256 3878
rect 24916 3806 24944 4012
rect 26112 3874 26140 4012
rect 27308 3942 27336 4012
rect 27296 3936 27348 3942
rect 27296 3878 27348 3884
rect 27712 3936 27764 3942
rect 27712 3878 27764 3884
rect 26100 3868 26152 3874
rect 26100 3810 26152 3816
rect 26516 3868 26568 3874
rect 26516 3810 26568 3816
rect 24904 3800 24956 3806
rect 24904 3742 24956 3748
rect 25320 3800 25372 3806
rect 25320 3742 25372 3748
rect 25332 480 25360 3742
rect 26528 480 26556 3810
rect 27724 480 27752 3878
rect 28412 3806 28440 4012
rect 29608 3874 29636 4012
rect 30712 3942 30740 4012
rect 30700 3936 30752 3942
rect 30700 3878 30752 3884
rect 29596 3868 29648 3874
rect 29596 3810 29648 3816
rect 30104 3868 30156 3874
rect 30104 3810 30156 3816
rect 28400 3800 28452 3806
rect 28400 3742 28452 3748
rect 28908 2848 28960 2854
rect 28908 2790 28960 2796
rect 28920 480 28948 2790
rect 30116 480 30144 3810
rect 31300 3800 31352 3806
rect 31908 3754 31936 4012
rect 32404 3936 32456 3942
rect 32404 3878 32456 3884
rect 31300 3742 31352 3748
rect 31312 480 31340 3742
rect 31864 3726 31936 3754
rect 31864 2854 31892 3726
rect 31852 2848 31904 2854
rect 31852 2790 31904 2796
rect 32416 480 32444 3878
rect 33104 3874 33132 4012
rect 33092 3868 33144 3874
rect 33092 3810 33144 3816
rect 33600 3868 33652 3874
rect 33600 3810 33652 3816
rect 33612 480 33640 3810
rect 34208 3806 34236 4012
rect 35404 3942 35432 4012
rect 35392 3936 35444 3942
rect 35392 3878 35444 3884
rect 36600 3874 36628 4012
rect 36588 3868 36640 3874
rect 36588 3810 36640 3816
rect 37188 3868 37240 3874
rect 37188 3810 37240 3816
rect 34196 3800 34248 3806
rect 34196 3742 34248 3748
rect 34796 3800 34848 3806
rect 34796 3742 34848 3748
rect 34808 480 34836 3742
rect 35992 2848 36044 2854
rect 35992 2790 36044 2796
rect 36004 480 36032 2790
rect 37200 480 37228 3810
rect 37704 3806 37732 4012
rect 38384 3936 38436 3942
rect 38384 3878 38436 3884
rect 37692 3800 37744 3806
rect 37692 3742 37744 3748
rect 38396 480 38424 3878
rect 38900 3754 38928 4012
rect 40004 3874 40032 4012
rect 41200 3942 41228 4012
rect 41188 3936 41240 3942
rect 41188 3878 41240 3884
rect 39992 3868 40044 3874
rect 39992 3810 40044 3816
rect 41880 3868 41932 3874
rect 41880 3810 41932 3816
rect 38856 3726 38928 3754
rect 40684 3800 40736 3806
rect 40684 3742 40736 3748
rect 38856 2854 38884 3726
rect 38844 2848 38896 2854
rect 38844 2790 38896 2796
rect 39580 2848 39632 2854
rect 39580 2790 39632 2796
rect 39592 480 39620 2790
rect 40696 480 40724 3742
rect 41892 480 41920 3810
rect 42396 3754 42424 4012
rect 43076 3936 43128 3942
rect 43076 3878 43128 3884
rect 42352 3726 42424 3754
rect 42352 2854 42380 3726
rect 42340 2848 42392 2854
rect 42340 2790 42392 2796
rect 43088 480 43116 3878
rect 43500 3806 43528 4012
rect 44696 3874 44724 4012
rect 45800 3942 45828 4012
rect 45788 3936 45840 3942
rect 45788 3878 45840 3884
rect 46664 3936 46716 3942
rect 46664 3878 46716 3884
rect 44684 3868 44736 3874
rect 44684 3810 44736 3816
rect 45468 3868 45520 3874
rect 45468 3810 45520 3816
rect 43488 3800 43540 3806
rect 43488 3742 43540 3748
rect 44272 3800 44324 3806
rect 44272 3742 44324 3748
rect 44284 480 44312 3742
rect 45480 480 45508 3810
rect 46676 480 46704 3878
rect 46996 3806 47024 4012
rect 48192 3874 48220 4012
rect 49296 3942 49324 4012
rect 49284 3936 49336 3942
rect 49284 3878 49336 3884
rect 50160 3936 50212 3942
rect 50160 3878 50212 3884
rect 48180 3868 48232 3874
rect 48180 3810 48232 3816
rect 48964 3868 49016 3874
rect 48964 3810 49016 3816
rect 46984 3800 47036 3806
rect 46984 3742 47036 3748
rect 47860 3800 47912 3806
rect 47860 3742 47912 3748
rect 47872 480 47900 3742
rect 48976 480 49004 3810
rect 50172 480 50200 3878
rect 50492 3806 50520 4012
rect 51596 3874 51624 4012
rect 52792 3942 52820 4012
rect 52780 3936 52832 3942
rect 52780 3878 52832 3884
rect 51584 3868 51636 3874
rect 51584 3810 51636 3816
rect 53748 3868 53800 3874
rect 53748 3810 53800 3816
rect 50480 3800 50532 3806
rect 50480 3742 50532 3748
rect 51356 3800 51408 3806
rect 51356 3742 51408 3748
rect 51368 480 51396 3742
rect 52552 740 52604 746
rect 52552 682 52604 688
rect 52564 480 52592 682
rect 53760 480 53788 3810
rect 53988 3806 54016 4012
rect 53976 3800 54028 3806
rect 53976 3742 54028 3748
rect 54944 3800 54996 3806
rect 55092 3754 55120 4012
rect 56048 3936 56100 3942
rect 56048 3878 56100 3884
rect 54944 3742 54996 3748
rect 54956 480 54984 3742
rect 55048 3726 55120 3754
rect 55048 746 55076 3726
rect 55036 740 55088 746
rect 55036 682 55088 688
rect 56060 480 56088 3878
rect 56288 3874 56316 4012
rect 56276 3868 56328 3874
rect 56276 3810 56328 3816
rect 57244 3868 57296 3874
rect 57244 3810 57296 3816
rect 57256 480 57284 3810
rect 57392 3806 57420 4012
rect 58588 3942 58616 4012
rect 58576 3936 58628 3942
rect 58576 3878 58628 3884
rect 59784 3874 59812 4012
rect 59772 3868 59824 3874
rect 59772 3810 59824 3816
rect 60888 3806 60916 4012
rect 62084 3890 62112 4012
rect 61948 3862 62112 3890
rect 57380 3800 57432 3806
rect 57380 3742 57432 3748
rect 58440 3800 58492 3806
rect 58440 3742 58492 3748
rect 60876 3800 60928 3806
rect 60876 3742 60928 3748
rect 58452 480 58480 3742
rect 60832 1352 60884 1358
rect 60832 1294 60884 1300
rect 59636 740 59688 746
rect 59636 682 59688 688
rect 59648 480 59676 682
rect 60844 480 60872 1294
rect 61948 746 61976 3862
rect 63280 3754 63308 4012
rect 64384 3890 64412 4012
rect 64384 3862 64460 3890
rect 64328 3800 64380 3806
rect 63280 3726 63356 3754
rect 64328 3742 64380 3748
rect 63224 3052 63276 3058
rect 63224 2994 63276 3000
rect 62028 2848 62080 2854
rect 62028 2790 62080 2796
rect 61936 740 61988 746
rect 61936 682 61988 688
rect 62040 480 62068 2790
rect 63236 480 63264 2994
rect 63328 1358 63356 3726
rect 63316 1352 63368 1358
rect 63316 1294 63368 1300
rect 64340 480 64368 3742
rect 64432 2854 64460 3862
rect 65580 3754 65608 4012
rect 66684 3806 66712 4012
rect 65536 3726 65608 3754
rect 66672 3800 66724 3806
rect 66672 3742 66724 3748
rect 67088 3800 67140 3806
rect 67880 3754 67908 4012
rect 69076 3806 69104 4012
rect 67088 3742 67140 3748
rect 65536 3058 65564 3726
rect 65524 3052 65576 3058
rect 65524 2994 65576 3000
rect 64420 2848 64472 2854
rect 64420 2790 64472 2796
rect 65524 2848 65576 2854
rect 65524 2790 65576 2796
rect 65536 480 65564 2790
rect 5234 326 5672 354
rect 5234 -960 5346 326
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 218 66802 480
rect 67100 218 67128 3742
rect 67836 3726 67908 3754
rect 69064 3800 69116 3806
rect 70180 3754 70208 4012
rect 69064 3742 69116 3748
rect 70136 3726 70208 3754
rect 70308 3800 70360 3806
rect 71376 3754 71404 4012
rect 71504 3868 71556 3874
rect 71504 3810 71556 3816
rect 70308 3742 70360 3748
rect 67836 2854 67864 3726
rect 67824 2848 67876 2854
rect 67824 2790 67876 2796
rect 70136 1358 70164 3726
rect 67916 1352 67968 1358
rect 67916 1294 67968 1300
rect 70124 1352 70176 1358
rect 70124 1294 70176 1300
rect 67928 480 67956 1294
rect 69112 604 69164 610
rect 69112 546 69164 552
rect 69124 480 69152 546
rect 70320 480 70348 3742
rect 71332 3726 71404 3754
rect 71332 610 71360 3726
rect 71320 604 71372 610
rect 71320 546 71372 552
rect 71516 480 71544 3810
rect 72480 3806 72508 4012
rect 72608 3936 72660 3942
rect 72608 3878 72660 3884
rect 72468 3800 72520 3806
rect 72468 3742 72520 3748
rect 72620 480 72648 3878
rect 73676 3874 73704 4012
rect 74872 3942 74900 4012
rect 74860 3936 74912 3942
rect 74860 3878 74912 3884
rect 73664 3868 73716 3874
rect 73664 3810 73716 3816
rect 75976 3806 76004 4012
rect 73804 3800 73856 3806
rect 73804 3742 73856 3748
rect 75964 3800 76016 3806
rect 77172 3754 77200 4012
rect 78276 3754 78304 4012
rect 78588 3868 78640 3874
rect 78588 3810 78640 3816
rect 75964 3742 76016 3748
rect 73816 480 73844 3742
rect 77128 3726 77200 3754
rect 78232 3726 78304 3754
rect 76196 1352 76248 1358
rect 76196 1294 76248 1300
rect 75000 1284 75052 1290
rect 75000 1226 75052 1232
rect 75012 480 75040 1226
rect 76208 480 76236 1294
rect 77128 1290 77156 3726
rect 78232 1358 78260 3726
rect 78220 1352 78272 1358
rect 78220 1294 78272 1300
rect 77116 1284 77168 1290
rect 77116 1226 77168 1232
rect 77392 1284 77444 1290
rect 77392 1226 77444 1232
rect 77404 480 77432 1226
rect 78600 480 78628 3810
rect 79472 3754 79500 4012
rect 80668 3874 80696 4012
rect 80656 3868 80708 3874
rect 80656 3810 80708 3816
rect 80888 3868 80940 3874
rect 80888 3810 80940 3816
rect 79428 3726 79500 3754
rect 79692 3800 79744 3806
rect 79692 3742 79744 3748
rect 79428 1290 79456 3726
rect 79416 1284 79468 1290
rect 79416 1226 79468 1232
rect 79704 480 79732 3742
rect 80900 480 80928 3810
rect 81772 3806 81800 4012
rect 82968 3874 82996 4012
rect 82956 3868 83008 3874
rect 82956 3810 83008 3816
rect 81760 3800 81812 3806
rect 84072 3754 84100 4012
rect 85268 3754 85296 4012
rect 86464 3754 86492 4012
rect 81760 3742 81812 3748
rect 84028 3726 84100 3754
rect 85224 3726 85296 3754
rect 86420 3726 86492 3754
rect 86868 3800 86920 3806
rect 87568 3754 87596 4012
rect 87972 3868 88024 3874
rect 87972 3810 88024 3816
rect 86868 3742 86920 3748
rect 83280 1352 83332 1358
rect 83280 1294 83332 1300
rect 82084 1284 82136 1290
rect 82084 1226 82136 1232
rect 82096 480 82124 1226
rect 83292 480 83320 1294
rect 84028 1290 84056 3726
rect 85224 1358 85252 3726
rect 85212 1352 85264 1358
rect 85212 1294 85264 1300
rect 85672 1352 85724 1358
rect 85672 1294 85724 1300
rect 84016 1284 84068 1290
rect 84016 1226 84068 1232
rect 84476 1284 84528 1290
rect 84476 1226 84528 1232
rect 84488 480 84516 1226
rect 85684 480 85712 1294
rect 86420 1290 86448 3726
rect 86408 1284 86460 1290
rect 86408 1226 86460 1232
rect 86880 480 86908 3742
rect 87524 3726 87596 3754
rect 87524 1358 87552 3726
rect 87512 1352 87564 1358
rect 87512 1294 87564 1300
rect 87984 480 88012 3810
rect 88764 3806 88792 4012
rect 89960 3874 89988 4012
rect 89948 3868 90000 3874
rect 89948 3810 90000 3816
rect 88752 3800 88804 3806
rect 91064 3754 91092 4012
rect 92260 3754 92288 4012
rect 93364 3754 93392 4012
rect 94560 3754 94588 4012
rect 88752 3742 88804 3748
rect 91020 3726 91092 3754
rect 92216 3726 92288 3754
rect 93320 3726 93392 3754
rect 94516 3726 94588 3754
rect 95148 3800 95200 3806
rect 95756 3754 95784 4012
rect 96252 3868 96304 3874
rect 96252 3810 96304 3816
rect 95148 3742 95200 3748
rect 91020 1358 91048 3726
rect 89168 1352 89220 1358
rect 89168 1294 89220 1300
rect 91008 1352 91060 1358
rect 91008 1294 91060 1300
rect 91560 1352 91612 1358
rect 91560 1294 91612 1300
rect 89180 480 89208 1294
rect 90364 1284 90416 1290
rect 90364 1226 90416 1232
rect 90376 480 90404 1226
rect 91572 480 91600 1294
rect 92216 1290 92244 3726
rect 93320 1358 93348 3726
rect 93308 1352 93360 1358
rect 93308 1294 93360 1300
rect 93952 1352 94004 1358
rect 93952 1294 94004 1300
rect 92204 1284 92256 1290
rect 92204 1226 92256 1232
rect 92756 1284 92808 1290
rect 92756 1226 92808 1232
rect 92768 480 92796 1226
rect 93964 480 93992 1294
rect 94516 1290 94544 3726
rect 94504 1284 94556 1290
rect 94504 1226 94556 1232
rect 95160 480 95188 3742
rect 95712 3726 95784 3754
rect 95712 1358 95740 3726
rect 95700 1352 95752 1358
rect 95700 1294 95752 1300
rect 96264 480 96292 3810
rect 96860 3806 96888 4012
rect 98056 3874 98084 4012
rect 98044 3868 98096 3874
rect 98044 3810 98096 3816
rect 96848 3800 96900 3806
rect 99160 3754 99188 4012
rect 100356 3754 100384 4012
rect 101552 3754 101580 4012
rect 102656 3754 102684 4012
rect 96848 3742 96900 3748
rect 99116 3726 99188 3754
rect 100312 3726 100384 3754
rect 101508 3726 101580 3754
rect 102612 3726 102684 3754
rect 103336 3800 103388 3806
rect 103852 3754 103880 4012
rect 104956 3806 104984 4012
rect 103336 3742 103388 3748
rect 99116 1358 99144 3726
rect 97448 1352 97500 1358
rect 97448 1294 97500 1300
rect 99104 1352 99156 1358
rect 99104 1294 99156 1300
rect 97460 480 97488 1294
rect 100312 1290 100340 3726
rect 101036 1352 101088 1358
rect 101036 1294 101088 1300
rect 98644 1284 98696 1290
rect 98644 1226 98696 1232
rect 100300 1284 100352 1290
rect 100300 1226 100352 1232
rect 98656 480 98684 1226
rect 99840 1216 99892 1222
rect 99840 1158 99892 1164
rect 99852 480 99880 1158
rect 101048 480 101076 1294
rect 101508 1222 101536 3726
rect 102612 1358 102640 3726
rect 102600 1352 102652 1358
rect 102600 1294 102652 1300
rect 102232 1284 102284 1290
rect 102232 1226 102284 1232
rect 101496 1216 101548 1222
rect 101496 1158 101548 1164
rect 102244 480 102272 1226
rect 103348 480 103376 3742
rect 103808 3726 103880 3754
rect 104944 3800 104996 3806
rect 106152 3754 106180 4012
rect 107348 3754 107376 4012
rect 108452 3754 108480 4012
rect 109648 3754 109676 4012
rect 110752 3754 110780 4012
rect 111948 3754 111976 4012
rect 113144 3754 113172 4012
rect 114248 3754 114276 4012
rect 115444 3754 115472 4012
rect 116640 3754 116668 4012
rect 117744 3754 117772 4012
rect 118940 3754 118968 4012
rect 120044 3754 120072 4012
rect 121240 3754 121268 4012
rect 122436 3754 122464 4012
rect 123540 3754 123568 4012
rect 104944 3742 104996 3748
rect 106108 3726 106180 3754
rect 107304 3726 107376 3754
rect 108408 3726 108480 3754
rect 109604 3726 109676 3754
rect 110708 3726 110780 3754
rect 111904 3726 111976 3754
rect 113100 3726 113172 3754
rect 114204 3726 114276 3754
rect 115400 3726 115472 3754
rect 116596 3726 116668 3754
rect 117700 3726 117772 3754
rect 118896 3726 118968 3754
rect 119264 3726 120072 3754
rect 121196 3726 121268 3754
rect 122392 3726 122464 3754
rect 123496 3726 123568 3754
rect 124736 3754 124764 4012
rect 125840 3754 125868 4012
rect 127036 3754 127064 4012
rect 128232 3754 128260 4012
rect 129336 3754 129364 4012
rect 130532 3754 130560 4012
rect 131636 3754 131664 4012
rect 132832 3754 132860 4012
rect 134028 3754 134056 4012
rect 135132 3754 135160 4012
rect 136328 3754 136356 4012
rect 137432 3754 137460 4012
rect 138628 3754 138656 4012
rect 139824 3754 139852 4012
rect 140928 3754 140956 4012
rect 142124 3754 142152 4012
rect 143320 3754 143348 4012
rect 144424 3754 144452 4012
rect 145620 3754 145648 4012
rect 146724 3754 146752 4012
rect 147920 3754 147948 4012
rect 149116 3754 149144 4012
rect 150220 3754 150248 4012
rect 151416 3754 151444 4012
rect 152520 3754 152548 4012
rect 153716 3754 153744 4012
rect 154912 3754 154940 4012
rect 156016 3754 156044 4012
rect 157212 3754 157240 4012
rect 158316 3754 158344 4012
rect 159512 3754 159540 4012
rect 160708 3754 160736 4012
rect 161812 3754 161840 4012
rect 163008 3754 163036 4012
rect 164112 3754 164140 4012
rect 165308 3754 165336 4012
rect 166504 3754 166532 4012
rect 167608 3754 167636 4012
rect 168804 3754 168832 4012
rect 170000 3754 170028 4012
rect 171104 3754 171132 4012
rect 172300 3754 172328 4012
rect 173404 3754 173432 4012
rect 174600 3754 174628 4012
rect 175796 3754 175824 4012
rect 176900 3754 176928 4012
rect 178096 3754 178124 4012
rect 179200 3754 179228 4012
rect 124736 3726 124812 3754
rect 103808 1290 103836 3726
rect 106108 1358 106136 3726
rect 104532 1352 104584 1358
rect 104532 1294 104584 1300
rect 106096 1352 106148 1358
rect 106096 1294 106148 1300
rect 106924 1352 106976 1358
rect 106924 1294 106976 1300
rect 103796 1284 103848 1290
rect 103796 1226 103848 1232
rect 104544 480 104572 1294
rect 105728 740 105780 746
rect 105728 682 105780 688
rect 105740 480 105768 682
rect 106936 480 106964 1294
rect 107304 746 107332 3726
rect 108408 1358 108436 3726
rect 108396 1352 108448 1358
rect 108396 1294 108448 1300
rect 109316 1352 109368 1358
rect 109316 1294 109368 1300
rect 108120 1284 108172 1290
rect 108120 1226 108172 1232
rect 107292 740 107344 746
rect 107292 682 107344 688
rect 108132 480 108160 1226
rect 109328 480 109356 1294
rect 109604 1290 109632 3726
rect 110708 1358 110736 3726
rect 110696 1352 110748 1358
rect 110696 1294 110748 1300
rect 111904 1290 111932 3726
rect 112812 1352 112864 1358
rect 112812 1294 112864 1300
rect 109592 1284 109644 1290
rect 109592 1226 109644 1232
rect 110512 1284 110564 1290
rect 110512 1226 110564 1232
rect 111892 1284 111944 1290
rect 111892 1226 111944 1232
rect 110524 480 110552 1226
rect 111616 1148 111668 1154
rect 111616 1090 111668 1096
rect 111628 480 111656 1090
rect 112824 480 112852 1294
rect 113100 1154 113128 3726
rect 114204 1358 114232 3726
rect 114192 1352 114244 1358
rect 114192 1294 114244 1300
rect 115204 1284 115256 1290
rect 115204 1226 115256 1232
rect 114008 1216 114060 1222
rect 114008 1158 114060 1164
rect 113088 1148 113140 1154
rect 113088 1090 113140 1096
rect 114020 480 114048 1158
rect 115216 480 115244 1226
rect 115400 1222 115428 3726
rect 116400 1352 116452 1358
rect 116400 1294 116452 1300
rect 115388 1216 115440 1222
rect 115388 1158 115440 1164
rect 116412 480 116440 1294
rect 116596 1290 116624 3726
rect 117700 1358 117728 3726
rect 117688 1352 117740 1358
rect 117688 1294 117740 1300
rect 118896 1290 118924 3726
rect 116584 1284 116636 1290
rect 116584 1226 116636 1232
rect 117596 1284 117648 1290
rect 117596 1226 117648 1232
rect 118884 1284 118936 1290
rect 118884 1226 118936 1232
rect 117608 480 117636 1226
rect 66690 190 67128 218
rect 66690 -960 66802 190
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 354 118874 480
rect 119264 354 119292 3726
rect 121196 1358 121224 3726
rect 119896 1352 119948 1358
rect 119896 1294 119948 1300
rect 121184 1352 121236 1358
rect 121184 1294 121236 1300
rect 119908 480 119936 1294
rect 122288 1284 122340 1290
rect 122288 1226 122340 1232
rect 121092 944 121144 950
rect 121092 886 121144 892
rect 121104 480 121132 886
rect 122300 480 122328 1226
rect 122392 950 122420 3726
rect 123496 1290 123524 3726
rect 123484 1284 123536 1290
rect 123484 1226 123536 1232
rect 124680 1284 124732 1290
rect 124680 1226 124732 1232
rect 123484 1148 123536 1154
rect 123484 1090 123536 1096
rect 122380 944 122432 950
rect 122380 886 122432 892
rect 123496 480 123524 1090
rect 124692 480 124720 1226
rect 124784 1154 124812 3726
rect 125796 3726 125868 3754
rect 126992 3726 127064 3754
rect 127176 3726 128260 3754
rect 129292 3726 129364 3754
rect 130488 3726 130560 3754
rect 131592 3726 131664 3754
rect 132788 3726 132860 3754
rect 133984 3726 134056 3754
rect 134168 3726 135160 3754
rect 135272 3726 136356 3754
rect 137388 3726 137460 3754
rect 138584 3726 138656 3754
rect 139780 3726 139852 3754
rect 140884 3726 140956 3754
rect 141712 3726 142152 3754
rect 142448 3726 143348 3754
rect 143552 3726 144452 3754
rect 145576 3726 145648 3754
rect 146680 3726 146752 3754
rect 147600 3726 147948 3754
rect 149072 3726 149144 3754
rect 149992 3726 150248 3754
rect 151096 3726 151444 3754
rect 151832 3726 152548 3754
rect 153488 3726 153744 3754
rect 154868 3726 154940 3754
rect 155880 3726 156044 3754
rect 156616 3726 157240 3754
rect 158272 3726 158344 3754
rect 159376 3726 159540 3754
rect 160112 3726 160736 3754
rect 161584 3726 161840 3754
rect 162964 3726 163036 3754
rect 164068 3726 164140 3754
rect 164896 3726 165336 3754
rect 166460 3726 166532 3754
rect 167564 3726 167636 3754
rect 168392 3726 168832 3754
rect 169956 3726 170028 3754
rect 170784 3726 171132 3754
rect 172256 3726 172328 3754
rect 173176 3726 173432 3754
rect 174280 3726 174628 3754
rect 175752 3726 175824 3754
rect 176672 3726 176928 3754
rect 178052 3726 178124 3754
rect 179064 3726 179228 3754
rect 180396 3754 180424 4012
rect 181592 3754 181620 4012
rect 182696 3754 182724 4012
rect 180396 3726 180472 3754
rect 125796 1290 125824 3726
rect 126992 1358 127020 3726
rect 125876 1352 125928 1358
rect 125876 1294 125928 1300
rect 126980 1352 127032 1358
rect 126980 1294 127032 1300
rect 125784 1284 125836 1290
rect 125784 1226 125836 1232
rect 124772 1148 124824 1154
rect 124772 1090 124824 1096
rect 125888 480 125916 1294
rect 127176 1170 127204 3726
rect 129292 1290 129320 3726
rect 130488 1358 130516 3726
rect 131592 1358 131620 3726
rect 132788 1358 132816 3726
rect 133984 1358 134012 3726
rect 129372 1352 129424 1358
rect 129372 1294 129424 1300
rect 130476 1352 130528 1358
rect 130476 1294 130528 1300
rect 130568 1352 130620 1358
rect 130568 1294 130620 1300
rect 131580 1352 131632 1358
rect 131580 1294 131632 1300
rect 131764 1352 131816 1358
rect 131764 1294 131816 1300
rect 132776 1352 132828 1358
rect 132776 1294 132828 1300
rect 132960 1352 133012 1358
rect 132960 1294 133012 1300
rect 133972 1352 134024 1358
rect 133972 1294 134024 1300
rect 128176 1284 128228 1290
rect 128176 1226 128228 1232
rect 129280 1284 129332 1290
rect 129280 1226 129332 1232
rect 126992 1142 127204 1170
rect 126992 480 127020 1142
rect 128188 480 128216 1226
rect 129384 480 129412 1294
rect 130580 480 130608 1294
rect 131776 480 131804 1294
rect 132972 480 133000 1294
rect 134168 480 134196 3726
rect 135272 480 135300 3726
rect 137388 1290 137416 3726
rect 138584 1358 138612 3726
rect 137652 1352 137704 1358
rect 137652 1294 137704 1300
rect 138572 1352 138624 1358
rect 138572 1294 138624 1300
rect 136456 1284 136508 1290
rect 136456 1226 136508 1232
rect 137376 1284 137428 1290
rect 137376 1226 137428 1232
rect 136468 480 136496 1226
rect 137664 480 137692 1294
rect 139780 1290 139808 3726
rect 140884 1290 140912 3726
rect 138848 1284 138900 1290
rect 138848 1226 138900 1232
rect 139768 1284 139820 1290
rect 139768 1226 139820 1232
rect 140044 1284 140096 1290
rect 140044 1226 140096 1232
rect 140872 1284 140924 1290
rect 140872 1226 140924 1232
rect 138860 480 138888 1226
rect 140056 480 140084 1226
rect 118762 326 119292 354
rect 118762 -960 118874 326
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 354 141322 480
rect 141712 354 141740 3726
rect 142448 480 142476 3726
rect 143552 480 143580 3726
rect 145576 1358 145604 3726
rect 146680 1358 146708 3726
rect 144736 1352 144788 1358
rect 144736 1294 144788 1300
rect 145564 1352 145616 1358
rect 145564 1294 145616 1300
rect 145932 1352 145984 1358
rect 145932 1294 145984 1300
rect 146668 1352 146720 1358
rect 146668 1294 146720 1300
rect 144748 480 144776 1294
rect 145944 480 145972 1294
rect 141210 326 141740 354
rect 141210 -960 141322 326
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 354 147210 480
rect 147600 354 147628 3726
rect 149072 1358 149100 3726
rect 148324 1352 148376 1358
rect 148324 1294 148376 1300
rect 149060 1352 149112 1358
rect 149060 1294 149112 1300
rect 148336 480 148364 1294
rect 147098 326 147628 354
rect 147098 -960 147210 326
rect 148294 -960 148406 480
rect 149490 354 149602 480
rect 149992 354 150020 3726
rect 149490 326 150020 354
rect 150594 354 150706 480
rect 151096 354 151124 3726
rect 151832 480 151860 3726
rect 150594 326 151124 354
rect 149490 -960 149602 326
rect 150594 -960 150706 326
rect 151790 -960 151902 480
rect 152986 354 153098 480
rect 153488 354 153516 3726
rect 154868 1358 154896 3726
rect 154212 1352 154264 1358
rect 154212 1294 154264 1300
rect 154856 1352 154908 1358
rect 154856 1294 154908 1300
rect 154224 480 154252 1294
rect 152986 326 153516 354
rect 152986 -960 153098 326
rect 154182 -960 154294 480
rect 155378 354 155490 480
rect 155880 354 155908 3726
rect 156616 480 156644 3726
rect 155378 326 155908 354
rect 155378 -960 155490 326
rect 156574 -960 156686 480
rect 157770 354 157882 480
rect 158272 354 158300 3726
rect 157770 326 158300 354
rect 158874 354 158986 480
rect 159376 354 159404 3726
rect 160112 480 160140 3726
rect 158874 326 159404 354
rect 157770 -960 157882 326
rect 158874 -960 158986 326
rect 160070 -960 160182 480
rect 161266 354 161378 480
rect 161584 354 161612 3726
rect 162964 1358 162992 3726
rect 162492 1352 162544 1358
rect 162492 1294 162544 1300
rect 162952 1352 163004 1358
rect 162952 1294 163004 1300
rect 162504 480 162532 1294
rect 161266 326 161612 354
rect 161266 -960 161378 326
rect 162462 -960 162574 480
rect 163658 354 163770 480
rect 164068 354 164096 3726
rect 164896 480 164924 3726
rect 163658 326 164096 354
rect 163658 -960 163770 326
rect 164854 -960 164966 480
rect 166050 354 166162 480
rect 166460 354 166488 3726
rect 166050 326 166488 354
rect 167154 354 167266 480
rect 167564 354 167592 3726
rect 168392 480 168420 3726
rect 167154 326 167592 354
rect 166050 -960 166162 326
rect 167154 -960 167266 326
rect 168350 -960 168462 480
rect 169546 354 169658 480
rect 169956 354 169984 3726
rect 170784 480 170812 3726
rect 169546 326 169984 354
rect 169546 -960 169658 326
rect 170742 -960 170854 480
rect 171938 354 172050 480
rect 172256 354 172284 3726
rect 173176 480 173204 3726
rect 174280 480 174308 3726
rect 171938 326 172284 354
rect 171938 -960 172050 326
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 354 175546 480
rect 175752 354 175780 3726
rect 176672 480 176700 3726
rect 175434 326 175780 354
rect 175434 -960 175546 326
rect 176630 -960 176742 480
rect 177826 354 177938 480
rect 178052 354 178080 3726
rect 179064 480 179092 3726
rect 177826 326 178080 354
rect 177826 -960 177938 326
rect 179022 -960 179134 480
rect 180218 218 180330 480
rect 180444 218 180472 3726
rect 181456 3726 181620 3754
rect 182560 3726 182724 3754
rect 183892 3754 183920 4012
rect 184996 3754 185024 4012
rect 186192 3754 186220 4012
rect 187388 3754 187416 4012
rect 183892 3726 183968 3754
rect 181456 480 181484 3726
rect 182560 480 182588 3726
rect 180218 190 180472 218
rect 180218 -960 180330 190
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 218 183826 480
rect 183940 218 183968 3726
rect 184952 3726 185024 3754
rect 186148 3726 186220 3754
rect 187344 3726 187416 3754
rect 188492 3754 188520 4012
rect 189688 3754 189716 4012
rect 190792 3754 190820 4012
rect 191988 3754 192016 4012
rect 193184 3754 193212 4012
rect 194288 3754 194316 4012
rect 195484 3754 195512 4012
rect 188492 3726 188568 3754
rect 189688 3726 189764 3754
rect 190792 3726 190868 3754
rect 191988 3726 192064 3754
rect 193184 3726 193260 3754
rect 194288 3726 194456 3754
rect 184952 480 184980 3726
rect 186148 480 186176 3726
rect 187344 480 187372 3726
rect 188540 480 188568 3726
rect 189736 480 189764 3726
rect 190840 480 190868 3726
rect 192036 480 192064 3726
rect 193232 480 193260 3726
rect 194428 480 194456 3726
rect 195440 3726 195512 3754
rect 196680 3754 196708 4012
rect 197784 3754 197812 4012
rect 198980 3754 199008 4012
rect 196680 3726 196848 3754
rect 197784 3726 197952 3754
rect 183714 190 183968 218
rect 183714 -960 183826 190
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195440 218 195468 3726
rect 196820 480 196848 3726
rect 197924 480 197952 3726
rect 198936 3726 199008 3754
rect 200084 3754 200112 4012
rect 201280 3754 201308 4012
rect 202476 3754 202504 4012
rect 203580 3754 203608 4012
rect 204776 3754 204804 4012
rect 205880 3754 205908 4012
rect 207076 3754 207104 4012
rect 208272 3754 208300 4012
rect 209376 3754 209404 4012
rect 210572 3754 210600 4012
rect 211676 3754 211704 4012
rect 212872 3754 212900 4012
rect 214068 3754 214096 4012
rect 215172 3754 215200 4012
rect 216368 3806 216396 4012
rect 216356 3800 216408 3806
rect 200084 3726 200344 3754
rect 201280 3726 201356 3754
rect 202476 3726 202736 3754
rect 203580 3726 203656 3754
rect 204776 3726 205128 3754
rect 205880 3726 206232 3754
rect 207076 3726 207152 3754
rect 208272 3726 208624 3754
rect 209376 3726 209728 3754
rect 210572 3726 211016 3754
rect 211676 3726 211752 3754
rect 212872 3726 213408 3754
rect 214068 3726 214512 3754
rect 215172 3726 215248 3754
rect 216356 3742 216408 3748
rect 216864 3800 216916 3806
rect 216864 3742 216916 3748
rect 217472 3754 217500 4012
rect 218668 3754 218696 4012
rect 219864 3754 219892 4012
rect 220968 3754 220996 4012
rect 222164 3806 222192 4012
rect 222152 3800 222204 3806
rect 195582 218 195694 480
rect 195440 190 195694 218
rect 195582 -960 195694 190
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198936 218 198964 3726
rect 200316 480 200344 3726
rect 199078 218 199190 480
rect 198936 190 199190 218
rect 199078 -960 199190 190
rect 200274 -960 200386 480
rect 201328 354 201356 3726
rect 202708 480 202736 3726
rect 201470 354 201582 480
rect 201328 326 201582 354
rect 201470 -960 201582 326
rect 202666 -960 202778 480
rect 203628 354 203656 3726
rect 205100 480 205128 3726
rect 206204 480 206232 3726
rect 203862 354 203974 480
rect 203628 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207124 354 207152 3726
rect 208596 480 208624 3726
rect 209700 626 209728 3726
rect 209700 598 209774 626
rect 209746 480 209774 598
rect 210988 480 211016 3726
rect 207358 354 207470 480
rect 207124 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209746 326 209862 480
rect 209750 -960 209862 326
rect 210946 -960 211058 480
rect 211724 354 211752 3726
rect 213380 480 213408 3726
rect 214484 480 214512 3726
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215220 354 215248 3726
rect 216876 480 216904 3742
rect 217472 3726 217640 3754
rect 218668 3726 219296 3754
rect 219864 3726 220032 3754
rect 220968 3726 221136 3754
rect 222152 3742 222204 3748
rect 222752 3800 222804 3806
rect 222752 3742 222804 3748
rect 223360 3754 223388 4012
rect 224464 3806 224492 4012
rect 224452 3800 224504 3806
rect 215638 354 215750 480
rect 215220 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 217612 354 217640 3726
rect 219268 480 219296 3726
rect 218030 354 218142 480
rect 217612 326 218142 354
rect 218030 -960 218142 326
rect 219226 -960 219338 480
rect 220004 354 220032 3726
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 3726
rect 222764 480 222792 3742
rect 223360 3726 223528 3754
rect 224452 3742 224504 3748
rect 225144 3800 225196 3806
rect 225144 3742 225196 3748
rect 225660 3754 225688 4012
rect 226764 3754 226792 4012
rect 227960 3754 227988 4012
rect 229156 3754 229184 4012
rect 230260 3806 230288 4012
rect 231456 3806 231484 4012
rect 232560 3806 232588 4012
rect 233756 3806 233784 4012
rect 230248 3800 230300 3806
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223500 354 223528 3726
rect 225156 480 225184 3742
rect 225660 3726 225920 3754
rect 226764 3726 227576 3754
rect 227960 3726 228312 3754
rect 229156 3726 229416 3754
rect 230248 3742 230300 3748
rect 231032 3800 231084 3806
rect 231032 3742 231084 3748
rect 231444 3800 231496 3806
rect 231444 3742 231496 3748
rect 232228 3800 232280 3806
rect 232228 3742 232280 3748
rect 232548 3800 232600 3806
rect 232548 3742 232600 3748
rect 233424 3800 233476 3806
rect 233424 3742 233476 3748
rect 233744 3800 233796 3806
rect 233744 3742 233796 3748
rect 234620 3800 234672 3806
rect 234620 3742 234672 3748
rect 234952 3754 234980 4012
rect 236056 3754 236084 4012
rect 237252 3806 237280 4012
rect 238356 3806 238384 4012
rect 239552 3806 239580 4012
rect 240748 3806 240776 4012
rect 241852 3806 241880 4012
rect 237240 3800 237292 3806
rect 223918 354 224030 480
rect 223500 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 225892 354 225920 3726
rect 227548 480 227576 3726
rect 226310 354 226422 480
rect 225892 326 226422 354
rect 226310 -960 226422 326
rect 227506 -960 227618 480
rect 228284 354 228312 3726
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 3726
rect 231044 480 231072 3742
rect 232240 480 232268 3742
rect 233436 480 233464 3742
rect 234632 480 234660 3742
rect 234952 3726 235856 3754
rect 236056 3726 236592 3754
rect 237240 3742 237292 3748
rect 238116 3800 238168 3806
rect 238116 3742 238168 3748
rect 238344 3800 238396 3806
rect 238344 3742 238396 3748
rect 239312 3800 239364 3806
rect 239312 3742 239364 3748
rect 239540 3800 239592 3806
rect 239540 3742 239592 3748
rect 240508 3800 240560 3806
rect 240508 3742 240560 3748
rect 240736 3800 240788 3806
rect 240736 3742 240788 3748
rect 241704 3800 241756 3806
rect 241704 3742 241756 3748
rect 241840 3800 241892 3806
rect 241840 3742 241892 3748
rect 242900 3800 242952 3806
rect 242900 3742 242952 3748
rect 243048 3754 243076 4012
rect 244152 3874 244180 4012
rect 244140 3868 244192 3874
rect 244140 3810 244192 3816
rect 245200 3868 245252 3874
rect 245200 3810 245252 3816
rect 235828 480 235856 3726
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 3726
rect 238128 480 238156 3742
rect 239324 480 239352 3742
rect 240520 480 240548 3742
rect 241716 480 241744 3742
rect 242912 480 242940 3742
rect 243048 3726 244136 3754
rect 244108 480 244136 3726
rect 245212 480 245240 3810
rect 245348 3806 245376 4012
rect 246544 3806 246572 4012
rect 247648 3942 247676 4012
rect 247636 3936 247688 3942
rect 247636 3878 247688 3884
rect 248604 3936 248656 3942
rect 248604 3878 248656 3884
rect 248844 3890 248872 4012
rect 245336 3800 245388 3806
rect 245336 3742 245388 3748
rect 246396 3800 246448 3806
rect 246396 3742 246448 3748
rect 246532 3800 246584 3806
rect 246532 3742 246584 3748
rect 247592 3800 247644 3806
rect 247592 3742 247644 3748
rect 246408 480 246436 3742
rect 247604 480 247632 3742
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 236982 -960 237094 326
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248616 354 248644 3878
rect 248844 3862 248920 3890
rect 248892 2854 248920 3862
rect 250040 3806 250068 4012
rect 251144 3890 251172 4012
rect 251100 3862 251172 3890
rect 250028 3800 250080 3806
rect 250028 3742 250080 3748
rect 251100 2854 251128 3862
rect 252340 3806 252368 4012
rect 253444 3890 253472 4012
rect 254640 3890 254668 4012
rect 253400 3862 253472 3890
rect 254596 3862 254668 3890
rect 251180 3800 251232 3806
rect 251180 3742 251232 3748
rect 252328 3800 252380 3806
rect 252328 3742 252380 3748
rect 248880 2848 248932 2854
rect 248880 2790 248932 2796
rect 249984 2848 250036 2854
rect 249984 2790 250036 2796
rect 251088 2848 251140 2854
rect 251088 2790 251140 2796
rect 249996 480 250024 2790
rect 251192 480 251220 3742
rect 253400 2922 253428 3862
rect 253480 3800 253532 3806
rect 253480 3742 253532 3748
rect 253388 2916 253440 2922
rect 253388 2858 253440 2864
rect 252376 2848 252428 2854
rect 252376 2790 252428 2796
rect 252388 480 252416 2790
rect 253492 480 253520 3742
rect 254596 2854 254624 3862
rect 255836 3806 255864 4012
rect 256940 3874 256968 4012
rect 256928 3868 256980 3874
rect 256928 3810 256980 3816
rect 258136 3806 258164 4012
rect 259240 3874 259268 4012
rect 258264 3868 258316 3874
rect 258264 3810 258316 3816
rect 259228 3868 259280 3874
rect 259228 3810 259280 3816
rect 255824 3800 255876 3806
rect 255824 3742 255876 3748
rect 257068 3800 257120 3806
rect 257068 3742 257120 3748
rect 258124 3800 258176 3806
rect 258124 3742 258176 3748
rect 254676 2916 254728 2922
rect 254676 2858 254728 2864
rect 254584 2848 254636 2854
rect 254584 2790 254636 2796
rect 254688 480 254716 2858
rect 255872 2848 255924 2854
rect 255872 2790 255924 2796
rect 255884 480 255912 2790
rect 257080 480 257108 3742
rect 258276 480 258304 3810
rect 260436 3806 260464 4012
rect 261632 3874 261660 4012
rect 260656 3868 260708 3874
rect 260656 3810 260708 3816
rect 261620 3868 261672 3874
rect 261620 3810 261672 3816
rect 259460 3800 259512 3806
rect 259460 3742 259512 3748
rect 260424 3800 260476 3806
rect 260424 3742 260476 3748
rect 259472 480 259500 3742
rect 260668 480 260696 3810
rect 262736 3806 262764 4012
rect 263932 3874 263960 4012
rect 262956 3868 263008 3874
rect 262956 3810 263008 3816
rect 263920 3868 263972 3874
rect 263920 3810 263972 3816
rect 261760 3800 261812 3806
rect 261760 3742 261812 3748
rect 262724 3800 262776 3806
rect 262724 3742 262776 3748
rect 261772 480 261800 3742
rect 262968 480 262996 3810
rect 265036 3806 265064 4012
rect 265348 3868 265400 3874
rect 265348 3810 265400 3816
rect 264152 3800 264204 3806
rect 264152 3742 264204 3748
rect 265024 3800 265076 3806
rect 265024 3742 265076 3748
rect 264164 480 264192 3742
rect 265360 480 265388 3810
rect 266232 3754 266260 4012
rect 267428 3806 267456 4012
rect 268532 3874 268560 4012
rect 268520 3868 268572 3874
rect 268520 3810 268572 3816
rect 269728 3806 269756 4012
rect 270832 3874 270860 4012
rect 270040 3868 270092 3874
rect 270040 3810 270092 3816
rect 270820 3868 270872 3874
rect 270820 3810 270872 3816
rect 266544 3800 266596 3806
rect 266232 3726 266308 3754
rect 266544 3742 266596 3748
rect 267416 3800 267468 3806
rect 267416 3742 267468 3748
rect 268844 3800 268896 3806
rect 268844 3742 268896 3748
rect 269716 3800 269768 3806
rect 269716 3742 269768 3748
rect 266280 1358 266308 3726
rect 266268 1352 266320 1358
rect 266268 1294 266320 1300
rect 266556 480 266584 3742
rect 267740 1352 267792 1358
rect 267740 1294 267792 1300
rect 267752 480 267780 1294
rect 268856 480 268884 3742
rect 270052 480 270080 3810
rect 272028 3806 272056 4012
rect 272432 3868 272484 3874
rect 272432 3810 272484 3816
rect 271236 3800 271288 3806
rect 271236 3742 271288 3748
rect 272016 3800 272068 3806
rect 272016 3742 272068 3748
rect 271248 480 271276 3742
rect 272444 480 272472 3810
rect 273224 3754 273252 4012
rect 273180 3726 273252 3754
rect 273628 3800 273680 3806
rect 273628 3742 273680 3748
rect 274328 3754 274356 4012
rect 275524 3874 275552 4012
rect 275512 3868 275564 3874
rect 275512 3810 275564 3816
rect 276720 3806 276748 4012
rect 277824 3874 277852 4012
rect 277124 3868 277176 3874
rect 277124 3810 277176 3816
rect 277812 3868 277864 3874
rect 277812 3810 277864 3816
rect 276708 3800 276760 3806
rect 273180 1358 273208 3726
rect 273168 1352 273220 1358
rect 273168 1294 273220 1300
rect 273640 480 273668 3742
rect 274328 3726 274404 3754
rect 276708 3742 276760 3748
rect 274376 746 274404 3726
rect 274824 1352 274876 1358
rect 274824 1294 274876 1300
rect 274364 740 274416 746
rect 274364 682 274416 688
rect 274836 480 274864 1294
rect 276020 740 276072 746
rect 276020 682 276072 688
rect 276032 480 276060 682
rect 277136 480 277164 3810
rect 279020 3806 279048 4012
rect 279516 3868 279568 3874
rect 279516 3810 279568 3816
rect 278320 3800 278372 3806
rect 278320 3742 278372 3748
rect 279008 3800 279060 3806
rect 279008 3742 279060 3748
rect 278332 480 278360 3742
rect 279528 480 279556 3810
rect 280124 3754 280152 4012
rect 280080 3726 280152 3754
rect 280712 3800 280764 3806
rect 280712 3742 280764 3748
rect 281320 3754 281348 4012
rect 282516 3754 282544 4012
rect 283620 3806 283648 4012
rect 284816 3874 284844 4012
rect 285920 3942 285948 4012
rect 285908 3936 285960 3942
rect 285908 3878 285960 3884
rect 284804 3868 284856 3874
rect 284804 3810 284856 3816
rect 286600 3868 286652 3874
rect 286600 3810 286652 3816
rect 283608 3800 283660 3806
rect 280080 1358 280108 3726
rect 280068 1352 280120 1358
rect 280068 1294 280120 1300
rect 280724 480 280752 3742
rect 281320 3726 281396 3754
rect 282516 3726 282592 3754
rect 283608 3742 283660 3748
rect 285404 3800 285456 3806
rect 285404 3742 285456 3748
rect 281368 1290 281396 3726
rect 282564 1358 282592 3726
rect 281908 1352 281960 1358
rect 281908 1294 281960 1300
rect 282552 1352 282604 1358
rect 282552 1294 282604 1300
rect 284300 1352 284352 1358
rect 284300 1294 284352 1300
rect 281356 1284 281408 1290
rect 281356 1226 281408 1232
rect 281920 480 281948 1294
rect 283104 1284 283156 1290
rect 283104 1226 283156 1232
rect 283116 480 283144 1226
rect 284312 480 284340 1294
rect 285416 480 285444 3742
rect 286612 480 286640 3810
rect 287116 3806 287144 4012
rect 287796 3936 287848 3942
rect 287796 3878 287848 3884
rect 287104 3800 287156 3806
rect 287104 3742 287156 3748
rect 287808 480 287836 3878
rect 288312 3754 288340 4012
rect 288992 3800 289044 3806
rect 288312 3726 288388 3754
rect 288992 3742 289044 3748
rect 289416 3754 289444 4012
rect 290612 3754 290640 4012
rect 291716 3806 291744 4012
rect 292912 3874 292940 4012
rect 292900 3868 292952 3874
rect 292900 3810 292952 3816
rect 294108 3806 294136 4012
rect 294880 3868 294932 3874
rect 294880 3810 294932 3816
rect 291704 3800 291756 3806
rect 288360 1358 288388 3726
rect 288348 1352 288400 1358
rect 288348 1294 288400 1300
rect 289004 480 289032 3742
rect 289416 3726 289492 3754
rect 290612 3726 290688 3754
rect 291704 3742 291756 3748
rect 293684 3800 293736 3806
rect 293684 3742 293736 3748
rect 294096 3800 294148 3806
rect 294096 3742 294148 3748
rect 289464 1290 289492 3726
rect 290188 1352 290240 1358
rect 290188 1294 290240 1300
rect 289452 1284 289504 1290
rect 289452 1226 289504 1232
rect 290200 480 290228 1294
rect 290660 610 290688 3726
rect 291384 1284 291436 1290
rect 291384 1226 291436 1232
rect 290648 604 290700 610
rect 290648 546 290700 552
rect 291396 480 291424 1226
rect 292580 604 292632 610
rect 292580 546 292632 552
rect 292592 480 292620 546
rect 293696 480 293724 3742
rect 294892 480 294920 3810
rect 295212 3754 295240 4012
rect 296076 3800 296128 3806
rect 295212 3726 295288 3754
rect 296076 3742 296128 3748
rect 296408 3754 296436 4012
rect 297512 3754 297540 4012
rect 298708 3806 298736 4012
rect 299904 3874 299932 4012
rect 299892 3868 299944 3874
rect 299892 3810 299944 3816
rect 301008 3806 301036 4012
rect 301964 3868 302016 3874
rect 301964 3810 302016 3816
rect 298696 3800 298748 3806
rect 295260 1358 295288 3726
rect 295248 1352 295300 1358
rect 295248 1294 295300 1300
rect 296088 480 296116 3742
rect 296408 3726 296484 3754
rect 297512 3726 297588 3754
rect 298696 3742 298748 3748
rect 300768 3800 300820 3806
rect 300768 3742 300820 3748
rect 300996 3800 301048 3806
rect 300996 3742 301048 3748
rect 296456 1290 296484 3726
rect 297560 1358 297588 3726
rect 297272 1352 297324 1358
rect 297272 1294 297324 1300
rect 297548 1352 297600 1358
rect 297548 1294 297600 1300
rect 299664 1352 299716 1358
rect 299664 1294 299716 1300
rect 296444 1284 296496 1290
rect 296444 1226 296496 1232
rect 297284 480 297312 1294
rect 298468 1284 298520 1290
rect 298468 1226 298520 1232
rect 298480 480 298508 1226
rect 299676 480 299704 1294
rect 300780 480 300808 3742
rect 301976 480 302004 3810
rect 302204 3754 302232 4012
rect 302160 3726 302232 3754
rect 303160 3800 303212 3806
rect 303160 3742 303212 3748
rect 303308 3754 303336 4012
rect 304504 3754 304532 4012
rect 305700 3754 305728 4012
rect 306804 3874 306832 4012
rect 306792 3868 306844 3874
rect 306792 3810 306844 3816
rect 308000 3806 308028 4012
rect 309048 3868 309100 3874
rect 309048 3810 309100 3816
rect 307988 3800 308040 3806
rect 302160 1358 302188 3726
rect 302148 1352 302200 1358
rect 302148 1294 302200 1300
rect 303172 480 303200 3742
rect 303308 3726 303384 3754
rect 304504 3726 304580 3754
rect 305700 3726 305776 3754
rect 307988 3742 308040 3748
rect 303356 1290 303384 3726
rect 304356 1352 304408 1358
rect 304356 1294 304408 1300
rect 303344 1284 303396 1290
rect 303344 1226 303396 1232
rect 304368 480 304396 1294
rect 304552 610 304580 3726
rect 305748 1358 305776 3726
rect 305736 1352 305788 1358
rect 305736 1294 305788 1300
rect 307944 1352 307996 1358
rect 307944 1294 307996 1300
rect 305552 1284 305604 1290
rect 305552 1226 305604 1232
rect 304540 604 304592 610
rect 304540 546 304592 552
rect 305564 480 305592 1226
rect 306748 604 306800 610
rect 306748 546 306800 552
rect 306760 480 306788 546
rect 307956 480 307984 1294
rect 309060 480 309088 3810
rect 309196 3754 309224 4012
rect 310300 3890 310328 4012
rect 311496 3890 311524 4012
rect 310300 3862 310376 3890
rect 311496 3862 311572 3890
rect 310244 3800 310296 3806
rect 309196 3726 309272 3754
rect 310244 3742 310296 3748
rect 309244 2854 309272 3726
rect 309232 2848 309284 2854
rect 309232 2790 309284 2796
rect 310256 480 310284 3742
rect 310348 1358 310376 3862
rect 311440 2848 311492 2854
rect 311440 2790 311492 2796
rect 310336 1352 310388 1358
rect 310336 1294 310388 1300
rect 311452 480 311480 2790
rect 311544 1222 311572 3862
rect 312600 3754 312628 4012
rect 312556 3726 312628 3754
rect 313796 3754 313824 4012
rect 314992 3754 315020 4012
rect 316096 3806 316124 4012
rect 316084 3800 316136 3806
rect 313796 3726 313872 3754
rect 314992 3726 315068 3754
rect 317292 3754 317320 4012
rect 316084 3742 316136 3748
rect 312556 1290 312584 3726
rect 313844 1358 313872 3726
rect 315040 2854 315068 3726
rect 317248 3726 317320 3754
rect 318396 3754 318424 4012
rect 318524 3800 318576 3806
rect 318396 3726 318472 3754
rect 318524 3742 318576 3748
rect 319592 3754 319620 4012
rect 320788 3754 320816 4012
rect 321892 3754 321920 4012
rect 323088 3806 323116 4012
rect 323076 3800 323128 3806
rect 315028 2848 315080 2854
rect 315028 2790 315080 2796
rect 317248 1358 317276 3726
rect 317328 2848 317380 2854
rect 317328 2790 317380 2796
rect 312636 1352 312688 1358
rect 312636 1294 312688 1300
rect 313832 1352 313884 1358
rect 313832 1294 313884 1300
rect 316224 1352 316276 1358
rect 316224 1294 316276 1300
rect 317236 1352 317288 1358
rect 317236 1294 317288 1300
rect 312544 1284 312596 1290
rect 312544 1226 312596 1232
rect 311532 1216 311584 1222
rect 311532 1158 311584 1164
rect 312648 480 312676 1294
rect 315028 1284 315080 1290
rect 315028 1226 315080 1232
rect 313832 1216 313884 1222
rect 313832 1158 313884 1164
rect 313844 480 313872 1158
rect 315040 480 315068 1226
rect 316236 480 316264 1294
rect 317340 480 317368 2790
rect 318444 1290 318472 3726
rect 318432 1284 318484 1290
rect 318432 1226 318484 1232
rect 318536 480 318564 3742
rect 319592 3726 319668 3754
rect 320788 3726 320864 3754
rect 321892 3726 321968 3754
rect 323076 3742 323128 3748
rect 324192 3754 324220 4012
rect 325388 3754 325416 4012
rect 325608 3800 325660 3806
rect 324192 3726 324268 3754
rect 325388 3726 325464 3754
rect 325608 3742 325660 3748
rect 326584 3754 326612 4012
rect 327688 3754 327716 4012
rect 328884 3754 328912 4012
rect 329988 3754 330016 4012
rect 331184 3754 331212 4012
rect 319640 1222 319668 3726
rect 319720 1352 319772 1358
rect 319720 1294 319772 1300
rect 319628 1216 319680 1222
rect 319628 1158 319680 1164
rect 319732 480 319760 1294
rect 320836 1154 320864 3726
rect 321940 1358 321968 3726
rect 321928 1352 321980 1358
rect 321928 1294 321980 1300
rect 320916 1284 320968 1290
rect 320916 1226 320968 1232
rect 320824 1148 320876 1154
rect 320824 1090 320876 1096
rect 320928 480 320956 1226
rect 322112 1216 322164 1222
rect 322112 1158 322164 1164
rect 322124 480 322152 1158
rect 323308 1148 323360 1154
rect 323308 1090 323360 1096
rect 323320 480 323348 1090
rect 324240 610 324268 3726
rect 325436 1358 325464 3726
rect 324412 1352 324464 1358
rect 324412 1294 324464 1300
rect 325424 1352 325476 1358
rect 325424 1294 325476 1300
rect 324228 604 324280 610
rect 324228 546 324280 552
rect 324424 480 324452 1294
rect 325620 480 325648 3742
rect 326584 3726 326660 3754
rect 327688 3726 327764 3754
rect 328884 3726 328960 3754
rect 329988 3726 330064 3754
rect 326632 1018 326660 3726
rect 327736 1222 327764 3726
rect 328932 1358 328960 3726
rect 328000 1352 328052 1358
rect 328000 1294 328052 1300
rect 328920 1352 328972 1358
rect 328920 1294 328972 1300
rect 327724 1216 327776 1222
rect 327724 1158 327776 1164
rect 326620 1012 326672 1018
rect 326620 954 326672 960
rect 326804 604 326856 610
rect 326804 546 326856 552
rect 326816 480 326844 546
rect 328012 480 328040 1294
rect 330036 1290 330064 3726
rect 331140 3726 331212 3754
rect 332380 3754 332408 4012
rect 333484 3754 333512 4012
rect 334680 3754 334708 4012
rect 335876 3754 335904 4012
rect 336980 3754 337008 4012
rect 338176 3754 338204 4012
rect 339280 3754 339308 4012
rect 340476 3754 340504 4012
rect 341672 3754 341700 4012
rect 342776 3754 342804 4012
rect 343972 3754 344000 4012
rect 345076 3754 345104 4012
rect 346272 3754 346300 4012
rect 347468 3754 347496 4012
rect 348572 3754 348600 4012
rect 349768 3754 349796 4012
rect 350872 3754 350900 4012
rect 352068 3754 352096 4012
rect 353264 3754 353292 4012
rect 332380 3726 332456 3754
rect 333484 3726 333560 3754
rect 334680 3726 334756 3754
rect 335876 3726 335952 3754
rect 336980 3726 337056 3754
rect 338176 3726 338252 3754
rect 339280 3726 339356 3754
rect 340476 3726 340552 3754
rect 341672 3726 341748 3754
rect 342776 3726 342852 3754
rect 343972 3726 344048 3754
rect 345076 3726 345152 3754
rect 346272 3726 346348 3754
rect 347468 3726 347544 3754
rect 348572 3726 348648 3754
rect 349768 3726 349844 3754
rect 350872 3726 350948 3754
rect 352068 3726 352144 3754
rect 330024 1284 330076 1290
rect 330024 1226 330076 1232
rect 331140 1222 331168 3726
rect 332428 1358 332456 3726
rect 331588 1352 331640 1358
rect 331588 1294 331640 1300
rect 332416 1352 332468 1358
rect 332416 1294 332468 1300
rect 330392 1216 330444 1222
rect 330392 1158 330444 1164
rect 331128 1216 331180 1222
rect 331128 1158 331180 1164
rect 329196 1012 329248 1018
rect 329196 954 329248 960
rect 329208 480 329236 954
rect 330404 480 330432 1158
rect 331600 480 331628 1294
rect 332692 1284 332744 1290
rect 332692 1226 332744 1232
rect 332704 480 332732 1226
rect 333532 746 333560 3726
rect 334728 1290 334756 3726
rect 335924 1358 335952 3726
rect 335084 1352 335136 1358
rect 335084 1294 335136 1300
rect 335912 1352 335964 1358
rect 335912 1294 335964 1300
rect 334716 1284 334768 1290
rect 334716 1226 334768 1232
rect 333888 1216 333940 1222
rect 333888 1158 333940 1164
rect 333520 740 333572 746
rect 333520 682 333572 688
rect 333900 480 333928 1158
rect 335096 480 335124 1294
rect 337028 1222 337056 3726
rect 337476 1284 337528 1290
rect 337476 1226 337528 1232
rect 337016 1216 337068 1222
rect 337016 1158 337068 1164
rect 336280 740 336332 746
rect 336280 682 336332 688
rect 336292 480 336320 682
rect 337488 480 337516 1226
rect 338224 746 338252 3726
rect 339328 1358 339356 3726
rect 338672 1352 338724 1358
rect 338672 1294 338724 1300
rect 339316 1352 339368 1358
rect 339316 1294 339368 1300
rect 338212 740 338264 746
rect 338212 682 338264 688
rect 338684 480 338712 1294
rect 340524 1290 340552 3726
rect 340512 1284 340564 1290
rect 340512 1226 340564 1232
rect 341720 1222 341748 3726
rect 342168 1352 342220 1358
rect 342168 1294 342220 1300
rect 339868 1216 339920 1222
rect 339868 1158 339920 1164
rect 341708 1216 341760 1222
rect 341708 1158 341760 1164
rect 339880 480 339908 1158
rect 340972 740 341024 746
rect 340972 682 341024 688
rect 340984 480 341012 682
rect 342180 480 342208 1294
rect 342824 746 342852 3726
rect 344020 1290 344048 3726
rect 345124 1358 345152 3726
rect 345112 1352 345164 1358
rect 345112 1294 345164 1300
rect 343364 1284 343416 1290
rect 343364 1226 343416 1232
rect 344008 1284 344060 1290
rect 344008 1226 344060 1232
rect 342812 740 342864 746
rect 342812 682 342864 688
rect 343376 480 343404 1226
rect 344560 1216 344612 1222
rect 344560 1158 344612 1164
rect 344572 480 344600 1158
rect 346320 746 346348 3726
rect 346952 1284 347004 1290
rect 346952 1226 347004 1232
rect 345756 740 345808 746
rect 345756 682 345808 688
rect 346308 740 346360 746
rect 346308 682 346360 688
rect 345768 480 345796 682
rect 346964 480 346992 1226
rect 347516 882 347544 3726
rect 348056 1352 348108 1358
rect 348056 1294 348108 1300
rect 347504 876 347556 882
rect 347504 818 347556 824
rect 348068 480 348096 1294
rect 348620 1290 348648 3726
rect 349816 1358 349844 3726
rect 349804 1352 349856 1358
rect 349804 1294 349856 1300
rect 348608 1284 348660 1290
rect 348608 1226 348660 1232
rect 350448 876 350500 882
rect 350448 818 350500 824
rect 349252 740 349304 746
rect 349252 682 349304 688
rect 349264 480 349292 682
rect 350460 480 350488 818
rect 350920 746 350948 3726
rect 352116 1290 352144 3726
rect 353220 3726 353292 3754
rect 354368 3754 354396 4012
rect 355564 3754 355592 4012
rect 356668 3754 356696 4012
rect 357864 3754 357892 4012
rect 359060 3754 359088 4012
rect 360164 3754 360192 4012
rect 354368 3726 354444 3754
rect 355564 3726 355640 3754
rect 356668 3726 356744 3754
rect 357864 3726 357940 3754
rect 359060 3726 359136 3754
rect 353220 1358 353248 3726
rect 352840 1352 352892 1358
rect 352840 1294 352892 1300
rect 353208 1352 353260 1358
rect 353208 1294 353260 1300
rect 351644 1284 351696 1290
rect 351644 1226 351696 1232
rect 352104 1284 352156 1290
rect 352104 1226 352156 1232
rect 350908 740 350960 746
rect 350908 682 350960 688
rect 351656 480 351684 1226
rect 352852 480 352880 1294
rect 354036 740 354088 746
rect 354036 682 354088 688
rect 354048 480 354076 682
rect 248758 354 248870 480
rect 248616 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 354416 66 354444 3726
rect 355612 1290 355640 3726
rect 356716 1358 356744 3726
rect 356336 1352 356388 1358
rect 356336 1294 356388 1300
rect 356704 1352 356756 1358
rect 356704 1294 356756 1300
rect 355232 1284 355284 1290
rect 355232 1226 355284 1232
rect 355600 1284 355652 1290
rect 355600 1226 355652 1232
rect 355244 480 355272 1226
rect 356348 480 356376 1294
rect 357912 1222 357940 3726
rect 359108 1290 359136 3726
rect 360120 3726 360192 3754
rect 361360 3754 361388 4012
rect 362556 3754 362584 4012
rect 363660 3754 363688 4012
rect 364856 3754 364884 4012
rect 365960 3754 365988 4012
rect 367156 3754 367184 4012
rect 368352 3754 368380 4012
rect 369456 3754 369484 4012
rect 370652 3754 370680 4012
rect 371756 3754 371784 4012
rect 372952 3754 372980 4012
rect 374148 3754 374176 4012
rect 375252 3754 375280 4012
rect 376448 3754 376476 4012
rect 361360 3726 361436 3754
rect 362556 3726 362632 3754
rect 363660 3726 363736 3754
rect 364856 3726 364932 3754
rect 365960 3726 366036 3754
rect 367156 3726 367232 3754
rect 368352 3726 368428 3754
rect 369456 3726 369532 3754
rect 370652 3726 370728 3754
rect 371756 3726 371832 3754
rect 372952 3726 373028 3754
rect 374148 3726 374224 3754
rect 375252 3726 375328 3754
rect 359924 1352 359976 1358
rect 359924 1294 359976 1300
rect 358728 1284 358780 1290
rect 358728 1226 358780 1232
rect 359096 1284 359148 1290
rect 359096 1226 359148 1232
rect 357900 1216 357952 1222
rect 357900 1158 357952 1164
rect 358740 480 358768 1226
rect 359936 480 359964 1294
rect 360120 1154 360148 3726
rect 361120 1216 361172 1222
rect 361120 1158 361172 1164
rect 360108 1148 360160 1154
rect 360108 1090 360160 1096
rect 361132 480 361160 1158
rect 361408 882 361436 3726
rect 362604 1358 362632 3726
rect 362592 1352 362644 1358
rect 362592 1294 362644 1300
rect 363708 1290 363736 3726
rect 362316 1284 362368 1290
rect 362316 1226 362368 1232
rect 363696 1284 363748 1290
rect 363696 1226 363748 1232
rect 361396 876 361448 882
rect 361396 818 361448 824
rect 362328 480 362356 1226
rect 364904 1222 364932 3726
rect 365812 1352 365864 1358
rect 365812 1294 365864 1300
rect 364892 1216 364944 1222
rect 364892 1158 364944 1164
rect 363512 1148 363564 1154
rect 363512 1090 363564 1096
rect 363524 480 363552 1090
rect 364616 876 364668 882
rect 364616 818 364668 824
rect 364628 480 364656 818
rect 365824 480 365852 1294
rect 366008 746 366036 3726
rect 367204 1358 367232 3726
rect 367192 1352 367244 1358
rect 367192 1294 367244 1300
rect 367008 1284 367060 1290
rect 367008 1226 367060 1232
rect 365996 740 366048 746
rect 365996 682 366048 688
rect 367020 480 367048 1226
rect 368204 1216 368256 1222
rect 368204 1158 368256 1164
rect 368216 480 368244 1158
rect 368400 882 368428 3726
rect 368388 876 368440 882
rect 368388 818 368440 824
rect 369504 746 369532 3726
rect 370700 1358 370728 3726
rect 370596 1352 370648 1358
rect 370596 1294 370648 1300
rect 370688 1352 370740 1358
rect 370688 1294 370740 1300
rect 369400 740 369452 746
rect 369400 682 369452 688
rect 369492 740 369544 746
rect 369492 682 369544 688
rect 369412 480 369440 682
rect 370608 480 370636 1294
rect 371804 882 371832 3726
rect 373000 1290 373028 3726
rect 374092 1352 374144 1358
rect 374092 1294 374144 1300
rect 372988 1284 373040 1290
rect 372988 1226 373040 1232
rect 371700 876 371752 882
rect 371700 818 371752 824
rect 371792 876 371844 882
rect 371792 818 371844 824
rect 371712 480 371740 818
rect 372896 740 372948 746
rect 372896 682 372948 688
rect 372908 480 372936 682
rect 374104 480 374132 1294
rect 374196 1018 374224 3726
rect 375300 1222 375328 3726
rect 376404 3726 376476 3754
rect 377552 3754 377580 4012
rect 378748 3754 378776 4012
rect 379944 3754 379972 4012
rect 377552 3726 377628 3754
rect 378748 3726 378824 3754
rect 376404 1358 376432 3726
rect 376392 1352 376444 1358
rect 376392 1294 376444 1300
rect 377600 1290 377628 3726
rect 376484 1284 376536 1290
rect 376484 1226 376536 1232
rect 377588 1284 377640 1290
rect 377588 1226 377640 1232
rect 375288 1216 375340 1222
rect 375288 1158 375340 1164
rect 374184 1012 374236 1018
rect 374184 954 374236 960
rect 375288 876 375340 882
rect 375288 818 375340 824
rect 375300 480 375328 818
rect 376496 480 376524 1226
rect 378796 1086 378824 3726
rect 379900 3726 379972 3754
rect 381048 3754 381076 4012
rect 382244 3754 382272 4012
rect 381048 3726 381124 3754
rect 378876 1216 378928 1222
rect 378876 1158 378928 1164
rect 378784 1080 378836 1086
rect 378784 1022 378836 1028
rect 377680 1012 377732 1018
rect 377680 954 377732 960
rect 377692 480 377720 954
rect 378888 480 378916 1158
rect 379900 1018 379928 3726
rect 379980 1352 380032 1358
rect 379980 1294 380032 1300
rect 379888 1012 379940 1018
rect 379888 954 379940 960
rect 379992 480 380020 1294
rect 381096 1222 381124 3726
rect 382200 3726 382272 3754
rect 383348 3754 383376 4012
rect 384544 3754 384572 4012
rect 385740 3754 385768 4012
rect 386844 3754 386872 4012
rect 388040 3754 388068 4012
rect 389236 3754 389264 4012
rect 390340 3754 390368 4012
rect 391536 3754 391564 4012
rect 392640 3754 392668 4012
rect 393836 3754 393864 4012
rect 395032 3754 395060 4012
rect 396136 3754 396164 4012
rect 397332 3754 397360 4012
rect 398436 3754 398464 4012
rect 399632 3754 399660 4012
rect 400828 3754 400856 4012
rect 401932 3754 401960 4012
rect 403128 3754 403156 4012
rect 404232 3754 404260 4012
rect 405428 3754 405456 4012
rect 406624 3754 406652 4012
rect 407728 3754 407756 4012
rect 408924 3754 408952 4012
rect 410028 3754 410056 4012
rect 411224 3754 411252 4012
rect 383348 3726 383424 3754
rect 384544 3726 384620 3754
rect 385740 3726 385816 3754
rect 386844 3726 386920 3754
rect 388040 3726 388116 3754
rect 389236 3726 389312 3754
rect 390340 3726 390416 3754
rect 391536 3726 391612 3754
rect 392640 3726 392716 3754
rect 393836 3726 393912 3754
rect 395032 3726 395108 3754
rect 396136 3726 396212 3754
rect 397332 3726 397408 3754
rect 398436 3726 398512 3754
rect 399632 3726 399708 3754
rect 400828 3726 400904 3754
rect 401932 3726 402008 3754
rect 403128 3726 403204 3754
rect 404232 3726 404308 3754
rect 405428 3726 405504 3754
rect 406624 3726 406700 3754
rect 407728 3726 407804 3754
rect 408924 3726 409000 3754
rect 410028 3726 410104 3754
rect 381176 1284 381228 1290
rect 381176 1226 381228 1232
rect 381084 1216 381136 1222
rect 381084 1158 381136 1164
rect 381188 480 381216 1226
rect 382200 1154 382228 3726
rect 382188 1148 382240 1154
rect 382188 1090 382240 1096
rect 382372 1080 382424 1086
rect 382372 1022 382424 1028
rect 382384 480 382412 1022
rect 354404 60 354456 66
rect 354404 2 354456 8
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 82 357614 480
rect 357360 66 357614 82
rect 357348 60 357614 66
rect 357400 54 357614 60
rect 357348 2 357400 8
rect 357502 -960 357614 54
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383396 134 383424 3726
rect 383568 1012 383620 1018
rect 383568 954 383620 960
rect 383580 480 383608 954
rect 384592 882 384620 3726
rect 385788 1358 385816 3726
rect 385776 1352 385828 1358
rect 385776 1294 385828 1300
rect 384764 1216 384816 1222
rect 384764 1158 384816 1164
rect 384580 876 384632 882
rect 384580 818 384632 824
rect 384776 480 384804 1158
rect 385960 1148 386012 1154
rect 385960 1090 386012 1096
rect 385972 480 386000 1090
rect 386892 1086 386920 3726
rect 388088 1290 388116 3726
rect 388076 1284 388128 1290
rect 388076 1226 388128 1232
rect 389284 1154 389312 3726
rect 389456 1352 389508 1358
rect 389456 1294 389508 1300
rect 389272 1148 389324 1154
rect 389272 1090 389324 1096
rect 386880 1080 386932 1086
rect 386880 1022 386932 1028
rect 388260 876 388312 882
rect 388260 818 388312 824
rect 388272 480 388300 818
rect 389468 480 389496 1294
rect 390388 1222 390416 3726
rect 390376 1216 390428 1222
rect 390376 1158 390428 1164
rect 390652 1080 390704 1086
rect 390652 1022 390704 1028
rect 390664 480 390692 1022
rect 391584 882 391612 3726
rect 391848 1284 391900 1290
rect 391848 1226 391900 1232
rect 391572 876 391624 882
rect 391572 818 391624 824
rect 391860 480 391888 1226
rect 383384 128 383436 134
rect 383384 70 383436 76
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 386788 128 386840 134
rect 387126 82 387238 480
rect 386840 76 387238 82
rect 386788 70 387238 76
rect 386800 54 387238 70
rect 387126 -960 387238 54
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392688 66 392716 3726
rect 393884 1290 393912 3726
rect 395080 1358 395108 3726
rect 395068 1352 395120 1358
rect 395068 1294 395120 1300
rect 393872 1284 393924 1290
rect 393872 1226 393924 1232
rect 396184 1222 396212 3726
rect 394240 1216 394292 1222
rect 394240 1158 394292 1164
rect 396172 1216 396224 1222
rect 396172 1158 396224 1164
rect 393044 1148 393096 1154
rect 393044 1090 393096 1096
rect 393056 480 393084 1090
rect 394252 480 394280 1158
rect 397380 882 397408 3726
rect 397736 1284 397788 1290
rect 397736 1226 397788 1232
rect 395344 876 395396 882
rect 395344 818 395396 824
rect 397368 876 397420 882
rect 397368 818 397420 824
rect 395356 480 395384 818
rect 397748 480 397776 1226
rect 398484 1154 398512 3726
rect 399680 1358 399708 3726
rect 398932 1352 398984 1358
rect 398932 1294 398984 1300
rect 399668 1352 399720 1358
rect 399668 1294 399720 1300
rect 398472 1148 398524 1154
rect 398472 1090 398524 1096
rect 398944 480 398972 1294
rect 400876 1222 400904 3726
rect 400128 1216 400180 1222
rect 400128 1158 400180 1164
rect 400864 1216 400916 1222
rect 400864 1158 400916 1164
rect 400140 480 400168 1158
rect 401324 876 401376 882
rect 401324 818 401376 824
rect 401336 480 401364 818
rect 392676 60 392728 66
rect 392676 2 392728 8
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 82 396622 480
rect 396184 66 396622 82
rect 396172 60 396622 66
rect 396224 54 396622 60
rect 396172 2 396224 8
rect 396510 -960 396622 54
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 401980 202 402008 3726
rect 403176 1290 403204 3726
rect 403624 1352 403676 1358
rect 403624 1294 403676 1300
rect 403164 1284 403216 1290
rect 403164 1226 403216 1232
rect 402520 1148 402572 1154
rect 402520 1090 402572 1096
rect 402532 480 402560 1090
rect 403636 480 403664 1294
rect 404280 1154 404308 3726
rect 405476 1358 405504 3726
rect 405464 1352 405516 1358
rect 405464 1294 405516 1300
rect 404820 1216 404872 1222
rect 404820 1158 404872 1164
rect 404268 1148 404320 1154
rect 404268 1090 404320 1096
rect 404832 480 404860 1158
rect 406672 882 406700 3726
rect 407212 1284 407264 1290
rect 407212 1226 407264 1232
rect 406660 876 406712 882
rect 406660 818 406712 824
rect 407224 480 407252 1226
rect 407776 1222 407804 3726
rect 407764 1216 407816 1222
rect 407764 1158 407816 1164
rect 408972 1154 409000 3726
rect 409604 1352 409656 1358
rect 409604 1294 409656 1300
rect 408408 1148 408460 1154
rect 408408 1090 408460 1096
rect 408960 1148 409012 1154
rect 408960 1090 409012 1096
rect 408420 480 408448 1090
rect 409616 480 409644 1294
rect 410076 1290 410104 3726
rect 411180 3726 411252 3754
rect 412420 3754 412448 4012
rect 413524 3754 413552 4012
rect 414720 3754 414748 4012
rect 415916 3754 415944 4012
rect 417020 3754 417048 4012
rect 418216 3754 418244 4012
rect 419320 3754 419348 4012
rect 420516 3754 420544 4012
rect 421712 3754 421740 4012
rect 422816 3754 422844 4012
rect 424012 3754 424040 4012
rect 425116 3754 425144 4012
rect 426312 3754 426340 4012
rect 427508 3754 427536 4012
rect 428612 3754 428640 4012
rect 429808 3754 429836 4012
rect 430912 3754 430940 4012
rect 432108 3754 432136 4012
rect 433304 3754 433332 4012
rect 434408 3754 434436 4012
rect 412420 3726 412496 3754
rect 413524 3726 413600 3754
rect 414720 3726 414796 3754
rect 415916 3726 415992 3754
rect 417020 3726 417096 3754
rect 418216 3726 418292 3754
rect 419320 3726 419396 3754
rect 420516 3726 420592 3754
rect 421712 3726 421788 3754
rect 422816 3726 422892 3754
rect 424012 3726 424088 3754
rect 425116 3726 425192 3754
rect 426312 3726 426388 3754
rect 427508 3726 427584 3754
rect 428612 3726 428688 3754
rect 429808 3726 429884 3754
rect 430912 3726 431080 3754
rect 432108 3726 432184 3754
rect 411180 2854 411208 3726
rect 411168 2848 411220 2854
rect 411168 2790 411220 2796
rect 410064 1284 410116 1290
rect 410064 1226 410116 1232
rect 411904 1216 411956 1222
rect 411904 1158 411956 1164
rect 410800 876 410852 882
rect 410800 818 410852 824
rect 410812 480 410840 818
rect 411916 480 411944 1158
rect 401968 196 402020 202
rect 401968 138 402020 144
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 218 406098 480
rect 405986 202 406240 218
rect 405986 196 406252 202
rect 405986 190 406200 196
rect 405986 -960 406098 190
rect 406200 138 406252 144
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412468 406 412496 3726
rect 413572 1358 413600 3726
rect 413560 1352 413612 1358
rect 413560 1294 413612 1300
rect 414296 1284 414348 1290
rect 414296 1226 414348 1232
rect 413100 1148 413152 1154
rect 413100 1090 413152 1096
rect 413112 480 413140 1090
rect 414308 480 414336 1226
rect 414768 1018 414796 3726
rect 415492 2848 415544 2854
rect 415492 2790 415544 2796
rect 414756 1012 414808 1018
rect 414756 954 414808 960
rect 415504 480 415532 2790
rect 415964 1154 415992 3726
rect 415952 1148 416004 1154
rect 415952 1090 416004 1096
rect 417068 1086 417096 3726
rect 417884 1352 417936 1358
rect 417884 1294 417936 1300
rect 417056 1080 417108 1086
rect 417056 1022 417108 1028
rect 416688 604 416740 610
rect 416688 546 416740 552
rect 416700 480 416728 546
rect 417896 480 417924 1294
rect 418264 1290 418292 3726
rect 418252 1284 418304 1290
rect 418252 1226 418304 1232
rect 418988 1012 419040 1018
rect 418988 954 419040 960
rect 419000 480 419028 954
rect 419368 882 419396 3726
rect 420564 1222 420592 3726
rect 420552 1216 420604 1222
rect 420552 1158 420604 1164
rect 420184 1148 420236 1154
rect 420184 1090 420236 1096
rect 419356 876 419408 882
rect 419356 818 419408 824
rect 420196 480 420224 1090
rect 421380 1080 421432 1086
rect 421380 1022 421432 1028
rect 421392 480 421420 1022
rect 412456 400 412508 406
rect 412456 342 412508 348
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 421760 134 421788 3726
rect 422864 1358 422892 3726
rect 422852 1352 422904 1358
rect 422852 1294 422904 1300
rect 422576 1284 422628 1290
rect 422576 1226 422628 1232
rect 422588 480 422616 1226
rect 424060 1018 424088 3726
rect 425164 1222 425192 3726
rect 426360 1290 426388 3726
rect 427556 1358 427584 3726
rect 427268 1352 427320 1358
rect 427268 1294 427320 1300
rect 427544 1352 427596 1358
rect 427544 1294 427596 1300
rect 426348 1284 426400 1290
rect 426348 1226 426400 1232
rect 424968 1216 425020 1222
rect 424968 1158 425020 1164
rect 425152 1216 425204 1222
rect 425152 1158 425204 1164
rect 424048 1012 424100 1018
rect 424048 954 424100 960
rect 423404 876 423456 882
rect 423404 818 423456 824
rect 421748 128 421800 134
rect 421748 70 421800 76
rect 422546 -960 422658 480
rect 423416 354 423444 818
rect 424980 480 425008 1158
rect 427280 480 427308 1294
rect 428660 1086 428688 3726
rect 429660 1216 429712 1222
rect 429660 1158 429712 1164
rect 428648 1080 428700 1086
rect 428648 1022 428700 1028
rect 428464 1012 428516 1018
rect 428464 954 428516 960
rect 428476 480 428504 954
rect 429672 480 429700 1158
rect 429856 1154 429884 3726
rect 430856 1284 430908 1290
rect 430856 1226 430908 1232
rect 429844 1148 429896 1154
rect 429844 1090 429896 1096
rect 430868 480 430896 1226
rect 423742 354 423854 480
rect 423416 326 423854 354
rect 423742 -960 423854 326
rect 424938 -960 425050 480
rect 425796 128 425848 134
rect 426134 82 426246 480
rect 425848 76 426246 82
rect 425796 70 426246 76
rect 425808 54 426246 70
rect 426134 -960 426246 54
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 431052 66 431080 3726
rect 431868 1352 431920 1358
rect 431868 1294 431920 1300
rect 431880 354 431908 1294
rect 432156 1018 432184 3726
rect 433260 3726 433332 3754
rect 434364 3726 434436 3754
rect 435604 3754 435632 4012
rect 436708 3754 436736 4012
rect 437904 3754 437932 4012
rect 439100 3754 439128 4012
rect 440204 3754 440232 4012
rect 435604 3726 435680 3754
rect 436708 3726 436784 3754
rect 437904 3726 437980 3754
rect 439100 3726 439176 3754
rect 433260 1358 433288 3726
rect 433248 1352 433300 1358
rect 433248 1294 433300 1300
rect 433248 1080 433300 1086
rect 433248 1022 433300 1028
rect 432144 1012 432196 1018
rect 432144 954 432196 960
rect 433260 480 433288 1022
rect 434364 882 434392 3726
rect 435652 1290 435680 3726
rect 435640 1284 435692 1290
rect 435640 1226 435692 1232
rect 436756 1154 436784 3726
rect 437848 1352 437900 1358
rect 437848 1294 437900 1300
rect 434444 1148 434496 1154
rect 434444 1090 434496 1096
rect 436744 1148 436796 1154
rect 436744 1090 436796 1096
rect 434352 876 434404 882
rect 434352 818 434404 824
rect 434456 480 434484 1090
rect 436744 1012 436796 1018
rect 436744 954 436796 960
rect 436756 480 436784 954
rect 437860 898 437888 1294
rect 437952 1086 437980 3726
rect 437940 1080 437992 1086
rect 437940 1022 437992 1028
rect 439148 1018 439176 3726
rect 440160 3726 440232 3754
rect 441400 3754 441428 4012
rect 442596 3754 442624 4012
rect 443700 3754 443728 4012
rect 444896 3754 444924 4012
rect 446000 3754 446028 4012
rect 447196 3754 447224 4012
rect 448392 3754 448420 4012
rect 449496 3754 449524 4012
rect 450692 3754 450720 4012
rect 451796 3754 451824 4012
rect 452992 3754 453020 4012
rect 454188 3754 454216 4012
rect 455292 3754 455320 4012
rect 456488 3754 456516 4012
rect 457592 3754 457620 4012
rect 458788 3754 458816 4012
rect 459984 3754 460012 4012
rect 461088 3754 461116 4012
rect 462284 3754 462312 4012
rect 441400 3726 441476 3754
rect 442596 3726 442672 3754
rect 443700 3726 443776 3754
rect 444896 3726 444972 3754
rect 446000 3726 446076 3754
rect 447196 3726 447272 3754
rect 448392 3726 448468 3754
rect 449496 3726 449572 3754
rect 450692 3726 450768 3754
rect 451796 3726 451872 3754
rect 452992 3726 453068 3754
rect 454188 3726 454264 3754
rect 455292 3726 455368 3754
rect 456488 3726 456564 3754
rect 457592 3726 457668 3754
rect 458788 3726 458864 3754
rect 459984 3726 460060 3754
rect 461088 3726 461164 3754
rect 440160 2854 440188 3726
rect 440148 2848 440200 2854
rect 440148 2790 440200 2796
rect 439964 1284 440016 1290
rect 439964 1226 440016 1232
rect 439136 1012 439188 1018
rect 439136 954 439188 960
rect 437860 870 437980 898
rect 437952 480 437980 870
rect 439136 876 439188 882
rect 439136 818 439188 824
rect 439148 480 439176 818
rect 432022 354 432134 480
rect 431880 326 432134 354
rect 431040 60 431092 66
rect 431040 2 431092 8
rect 432022 -960 432134 326
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 82 435630 480
rect 435192 66 435630 82
rect 435180 60 435630 66
rect 435232 54 435630 60
rect 435180 2 435232 8
rect 435518 -960 435630 54
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 439976 354 440004 1226
rect 441448 1222 441476 3726
rect 442644 1358 442672 3726
rect 442632 1352 442684 1358
rect 442632 1294 442684 1300
rect 443748 1290 443776 3726
rect 443736 1284 443788 1290
rect 443736 1226 443788 1232
rect 441436 1216 441488 1222
rect 441436 1158 441488 1164
rect 441528 1148 441580 1154
rect 441528 1090 441580 1096
rect 441540 480 441568 1090
rect 442632 1080 442684 1086
rect 442632 1022 442684 1028
rect 442644 480 442672 1022
rect 443828 1012 443880 1018
rect 443828 954 443880 960
rect 443840 480 443868 954
rect 444944 882 444972 3726
rect 445024 2848 445076 2854
rect 445024 2790 445076 2796
rect 444932 876 444984 882
rect 444932 818 444984 824
rect 445036 480 445064 2790
rect 445852 1216 445904 1222
rect 445852 1158 445904 1164
rect 440302 354 440414 480
rect 439976 326 440414 354
rect 440302 -960 440414 326
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445864 354 445892 1158
rect 446048 1154 446076 3726
rect 447244 1222 447272 3726
rect 448440 1358 448468 3726
rect 449544 2854 449572 3726
rect 449532 2848 449584 2854
rect 449532 2790 449584 2796
rect 447416 1352 447468 1358
rect 447416 1294 447468 1300
rect 448428 1352 448480 1358
rect 448428 1294 448480 1300
rect 447232 1216 447284 1222
rect 447232 1158 447284 1164
rect 446036 1148 446088 1154
rect 446036 1090 446088 1096
rect 447428 480 447456 1294
rect 450740 1290 450768 3726
rect 448244 1284 448296 1290
rect 448244 1226 448296 1232
rect 450728 1284 450780 1290
rect 450728 1226 450780 1232
rect 446190 354 446302 480
rect 445864 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448256 354 448284 1226
rect 450912 1148 450964 1154
rect 450912 1090 450964 1096
rect 449808 876 449860 882
rect 449808 818 449860 824
rect 449820 480 449848 818
rect 450924 480 450952 1090
rect 451844 746 451872 3726
rect 452108 1216 452160 1222
rect 452108 1158 452160 1164
rect 451832 740 451884 746
rect 451832 682 451884 688
rect 452120 480 452148 1158
rect 453040 1018 453068 3726
rect 453304 1352 453356 1358
rect 453304 1294 453356 1300
rect 453028 1012 453080 1018
rect 453028 954 453080 960
rect 453316 480 453344 1294
rect 454236 1222 454264 3726
rect 454500 2848 454552 2854
rect 454500 2790 454552 2796
rect 454224 1216 454276 1222
rect 454224 1158 454276 1164
rect 454512 480 454540 2790
rect 455340 1086 455368 3726
rect 456536 1290 456564 3726
rect 455696 1284 455748 1290
rect 455696 1226 455748 1232
rect 456524 1284 456576 1290
rect 456524 1226 456576 1232
rect 455328 1080 455380 1086
rect 455328 1022 455380 1028
rect 455708 480 455736 1226
rect 457640 1154 457668 3726
rect 458836 1358 458864 3726
rect 458824 1352 458876 1358
rect 458824 1294 458876 1300
rect 460032 1222 460060 3726
rect 459192 1216 459244 1222
rect 459192 1158 459244 1164
rect 460020 1216 460072 1222
rect 460020 1158 460072 1164
rect 457628 1148 457680 1154
rect 457628 1090 457680 1096
rect 458088 1012 458140 1018
rect 458088 954 458140 960
rect 456524 740 456576 746
rect 456524 682 456576 688
rect 448582 354 448694 480
rect 448256 326 448694 354
rect 448582 -960 448694 326
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456536 354 456564 682
rect 458100 480 458128 954
rect 459204 480 459232 1158
rect 460020 1080 460072 1086
rect 460020 1022 460072 1028
rect 456862 354 456974 480
rect 456536 326 456974 354
rect 456862 -960 456974 326
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460032 354 460060 1022
rect 461136 882 461164 3726
rect 462240 3726 462312 3754
rect 463388 3754 463416 4012
rect 464584 3754 464612 4012
rect 465780 3754 465808 4012
rect 466884 3754 466912 4012
rect 468080 3754 468108 4012
rect 469276 3754 469304 4012
rect 470380 3754 470408 4012
rect 471576 3754 471604 4012
rect 472680 3754 472708 4012
rect 473876 3754 473904 4012
rect 475072 3754 475100 4012
rect 476176 3754 476204 4012
rect 477372 3754 477400 4012
rect 478476 3754 478504 4012
rect 479672 3754 479700 4012
rect 480868 3754 480896 4012
rect 481972 3754 482000 4012
rect 483168 3754 483196 4012
rect 484272 3754 484300 4012
rect 485468 3754 485496 4012
rect 486664 3754 486692 4012
rect 487768 3754 487796 4012
rect 488964 3754 488992 4012
rect 490068 3754 490096 4012
rect 491264 3754 491292 4012
rect 463388 3726 463464 3754
rect 464584 3726 464660 3754
rect 465780 3726 465856 3754
rect 466884 3726 466960 3754
rect 468080 3726 468156 3754
rect 469276 3726 469352 3754
rect 470380 3726 470456 3754
rect 471576 3726 471652 3754
rect 472680 3726 472756 3754
rect 473876 3726 473952 3754
rect 475072 3726 475148 3754
rect 476176 3726 476252 3754
rect 477372 3726 477448 3754
rect 478476 3726 478552 3754
rect 479672 3726 479748 3754
rect 480868 3726 480944 3754
rect 481972 3726 482048 3754
rect 483168 3726 483244 3754
rect 484272 3726 484348 3754
rect 485468 3726 485544 3754
rect 486664 3726 486740 3754
rect 487768 3726 487844 3754
rect 488964 3726 489040 3754
rect 490068 3726 490144 3754
rect 462240 1290 462268 3726
rect 461584 1284 461636 1290
rect 461584 1226 461636 1232
rect 462228 1284 462280 1290
rect 462228 1226 462280 1232
rect 461124 876 461176 882
rect 461124 818 461176 824
rect 461596 480 461624 1226
rect 462412 1148 462464 1154
rect 462412 1090 462464 1096
rect 460358 354 460470 480
rect 460032 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462424 354 462452 1090
rect 463436 950 463464 3726
rect 463976 1352 464028 1358
rect 463976 1294 464028 1300
rect 463424 944 463476 950
rect 463424 886 463476 892
rect 463988 480 464016 1294
rect 464632 1154 464660 3726
rect 464804 1216 464856 1222
rect 464804 1158 464856 1164
rect 464620 1148 464672 1154
rect 464620 1090 464672 1096
rect 462750 354 462862 480
rect 462424 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 464816 354 464844 1158
rect 465828 1086 465856 3726
rect 465816 1080 465868 1086
rect 465816 1022 465868 1028
rect 466932 1018 466960 3726
rect 468128 1358 468156 3726
rect 468116 1352 468168 1358
rect 468116 1294 468168 1300
rect 467472 1284 467524 1290
rect 467472 1226 467524 1232
rect 466920 1012 466972 1018
rect 466920 954 466972 960
rect 466276 876 466328 882
rect 466276 818 466328 824
rect 466288 480 466316 818
rect 467484 480 467512 1226
rect 468300 944 468352 950
rect 468300 886 468352 892
rect 465142 354 465254 480
rect 464816 326 465254 354
rect 465142 -960 465254 326
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468312 354 468340 886
rect 468638 354 468750 480
rect 468312 326 468750 354
rect 468638 -960 468750 326
rect 469324 66 469352 3726
rect 470428 1222 470456 3726
rect 471624 1290 471652 3726
rect 471612 1284 471664 1290
rect 471612 1226 471664 1232
rect 470416 1216 470468 1222
rect 470416 1158 470468 1164
rect 472728 1154 472756 3726
rect 473084 1352 473136 1358
rect 473084 1294 473136 1300
rect 469864 1148 469916 1154
rect 469864 1090 469916 1096
rect 472716 1148 472768 1154
rect 472716 1090 472768 1096
rect 469876 480 469904 1090
rect 470692 1080 470744 1086
rect 470692 1022 470744 1028
rect 469312 60 469364 66
rect 469312 2 469364 8
rect 469834 -960 469946 480
rect 470704 354 470732 1022
rect 472256 1012 472308 1018
rect 472256 954 472308 960
rect 472268 480 472296 954
rect 471030 354 471142 480
rect 470704 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473096 354 473124 1294
rect 473924 1086 473952 3726
rect 475120 1358 475148 3726
rect 475108 1352 475160 1358
rect 475108 1294 475160 1300
rect 475752 1216 475804 1222
rect 475752 1158 475804 1164
rect 473912 1080 473964 1086
rect 473912 1022 473964 1028
rect 475764 480 475792 1158
rect 476224 1018 476252 3726
rect 476580 1284 476632 1290
rect 476580 1226 476632 1232
rect 476212 1012 476264 1018
rect 476212 954 476264 960
rect 473422 354 473534 480
rect 473096 326 473534 354
rect 473422 -960 473534 326
rect 474526 82 474638 480
rect 474200 66 474638 82
rect 474188 60 474638 66
rect 474240 54 474638 60
rect 474188 2 474240 8
rect 474526 -960 474638 54
rect 475722 -960 475834 480
rect 476592 354 476620 1226
rect 477420 1222 477448 3726
rect 478524 2854 478552 3726
rect 478512 2848 478564 2854
rect 478512 2790 478564 2796
rect 477408 1216 477460 1222
rect 477408 1158 477460 1164
rect 478144 1148 478196 1154
rect 478144 1090 478196 1096
rect 478156 480 478184 1090
rect 478972 1080 479024 1086
rect 478972 1022 479024 1028
rect 476918 354 477030 480
rect 476592 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 478984 354 479012 1022
rect 479720 950 479748 3726
rect 480536 1352 480588 1358
rect 480536 1294 480588 1300
rect 479708 944 479760 950
rect 479708 886 479760 892
rect 480548 480 480576 1294
rect 480916 1290 480944 3726
rect 480904 1284 480956 1290
rect 480904 1226 480956 1232
rect 482020 1086 482048 3726
rect 483216 1222 483244 3726
rect 484032 2848 484084 2854
rect 484032 2790 484084 2796
rect 482468 1216 482520 1222
rect 482468 1158 482520 1164
rect 483204 1216 483256 1222
rect 483204 1158 483256 1164
rect 482008 1080 482060 1086
rect 482008 1022 482060 1028
rect 481364 1012 481416 1018
rect 481364 954 481416 960
rect 479310 354 479422 480
rect 478984 326 479422 354
rect 479310 -960 479422 326
rect 480506 -960 480618 480
rect 481376 354 481404 954
rect 481702 354 481814 480
rect 481376 326 481814 354
rect 482480 354 482508 1158
rect 484044 480 484072 2790
rect 484320 882 484348 3726
rect 485516 1358 485544 3726
rect 485504 1352 485556 1358
rect 485504 1294 485556 1300
rect 486424 1284 486476 1290
rect 486424 1226 486476 1232
rect 484860 944 484912 950
rect 484860 886 484912 892
rect 484308 876 484360 882
rect 484308 818 484360 824
rect 482806 354 482918 480
rect 482480 326 482918 354
rect 481702 -960 481814 326
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484872 354 484900 886
rect 486436 480 486464 1226
rect 486712 1154 486740 3726
rect 487816 2854 487844 3726
rect 487804 2848 487856 2854
rect 487804 2790 487856 2796
rect 488816 1216 488868 1222
rect 488816 1158 488868 1164
rect 486700 1148 486752 1154
rect 486700 1090 486752 1096
rect 487252 1080 487304 1086
rect 487252 1022 487304 1028
rect 485198 354 485310 480
rect 484872 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487264 354 487292 1022
rect 488828 480 488856 1158
rect 489012 1018 489040 3726
rect 490116 1222 490144 3726
rect 491220 3726 491292 3754
rect 492460 3754 492488 4012
rect 493564 3754 493592 4012
rect 494760 3754 494788 4012
rect 495956 3754 495984 4012
rect 497060 3754 497088 4012
rect 498256 3754 498284 4012
rect 499360 3754 499388 4012
rect 500556 3754 500584 4012
rect 501752 3754 501780 4012
rect 502856 3754 502884 4012
rect 504052 3754 504080 4012
rect 505156 3754 505184 4012
rect 506352 3754 506380 4012
rect 507548 3754 507576 4012
rect 508652 3754 508680 4012
rect 509848 3754 509876 4012
rect 510952 3754 510980 4012
rect 512148 3754 512176 4012
rect 513344 3754 513372 4012
rect 492460 3726 492536 3754
rect 493564 3726 493640 3754
rect 494760 3726 494836 3754
rect 495956 3726 496032 3754
rect 497060 3726 497136 3754
rect 498256 3726 498332 3754
rect 499360 3726 499436 3754
rect 500556 3726 500632 3754
rect 501752 3726 501828 3754
rect 502856 3726 502932 3754
rect 504052 3726 504128 3754
rect 505156 3726 505232 3754
rect 506352 3726 506428 3754
rect 507548 3726 507624 3754
rect 508652 3726 508728 3754
rect 509848 3726 509924 3754
rect 510952 3726 511028 3754
rect 512148 3726 512224 3754
rect 490748 1352 490800 1358
rect 490748 1294 490800 1300
rect 490104 1216 490156 1222
rect 490104 1158 490156 1164
rect 489000 1012 489052 1018
rect 489000 954 489052 960
rect 489920 876 489972 882
rect 489920 818 489972 824
rect 489932 480 489960 818
rect 487590 354 487702 480
rect 487264 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 1294
rect 491220 1086 491248 3726
rect 492508 1290 492536 3726
rect 493508 2848 493560 2854
rect 493508 2790 493560 2796
rect 492496 1284 492548 1290
rect 492496 1226 492548 1232
rect 492312 1148 492364 1154
rect 492312 1090 492364 1096
rect 491208 1080 491260 1086
rect 491208 1022 491260 1028
rect 492324 480 492352 1090
rect 493520 480 493548 2790
rect 493612 950 493640 3726
rect 494808 1018 494836 3726
rect 495532 1216 495584 1222
rect 495532 1158 495584 1164
rect 494704 1012 494756 1018
rect 494704 954 494756 960
rect 494796 1012 494848 1018
rect 494796 954 494848 960
rect 493600 944 493652 950
rect 493600 886 493652 892
rect 494716 480 494744 954
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495544 354 495572 1158
rect 496004 882 496032 3726
rect 497108 1358 497136 3726
rect 497096 1352 497148 1358
rect 497096 1294 497148 1300
rect 498304 1290 498332 3726
rect 498200 1284 498252 1290
rect 498200 1226 498252 1232
rect 498292 1284 498344 1290
rect 498292 1226 498344 1232
rect 497096 1080 497148 1086
rect 497096 1022 497148 1028
rect 495992 876 496044 882
rect 495992 818 496044 824
rect 497108 480 497136 1022
rect 498212 480 498240 1226
rect 499408 1086 499436 3726
rect 500604 1154 500632 3726
rect 500592 1148 500644 1154
rect 500592 1090 500644 1096
rect 499396 1080 499448 1086
rect 499396 1022 499448 1028
rect 501800 1018 501828 3726
rect 500592 1012 500644 1018
rect 500592 954 500644 960
rect 501788 1012 501840 1018
rect 501788 954 501840 960
rect 499396 944 499448 950
rect 499396 886 499448 892
rect 499408 480 499436 886
rect 500604 480 500632 954
rect 502904 950 502932 3726
rect 504100 1358 504128 3726
rect 502984 1352 503036 1358
rect 502984 1294 503036 1300
rect 504088 1352 504140 1358
rect 504088 1294 504140 1300
rect 502892 944 502944 950
rect 502892 886 502944 892
rect 501788 876 501840 882
rect 501788 818 501840 824
rect 501800 480 501828 818
rect 502996 480 503024 1294
rect 503812 1284 503864 1290
rect 503812 1226 503864 1232
rect 495870 354 495982 480
rect 495544 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503824 354 503852 1226
rect 505204 1222 505232 3726
rect 506400 2922 506428 3726
rect 506388 2916 506440 2922
rect 506388 2858 506440 2864
rect 507596 2854 507624 3726
rect 507584 2848 507636 2854
rect 507584 2790 507636 2796
rect 505192 1216 505244 1222
rect 505192 1158 505244 1164
rect 506480 1148 506532 1154
rect 506480 1090 506532 1096
rect 505376 1080 505428 1086
rect 505376 1022 505428 1028
rect 505388 480 505416 1022
rect 506492 480 506520 1090
rect 508700 1086 508728 3726
rect 509700 1352 509752 1358
rect 509700 1294 509752 1300
rect 508688 1080 508740 1086
rect 508688 1022 508740 1028
rect 507308 1012 507360 1018
rect 507308 954 507360 960
rect 504150 354 504262 480
rect 503824 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507320 354 507348 954
rect 508872 944 508924 950
rect 508872 886 508924 892
rect 508884 480 508912 886
rect 507646 354 507758 480
rect 507320 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509712 354 509740 1294
rect 509896 1290 509924 3726
rect 509884 1284 509936 1290
rect 509884 1226 509936 1232
rect 511000 1154 511028 3726
rect 511264 1216 511316 1222
rect 511264 1158 511316 1164
rect 510988 1148 511040 1154
rect 510988 1090 511040 1096
rect 511276 480 511304 1158
rect 512196 1018 512224 3726
rect 513300 3726 513372 3754
rect 514448 3754 514476 4012
rect 515644 3754 515672 4012
rect 516748 3754 516776 4012
rect 517944 3754 517972 4012
rect 519140 3754 519168 4012
rect 520244 3754 520272 4012
rect 514448 3726 514524 3754
rect 515644 3726 515720 3754
rect 516748 3726 516824 3754
rect 517944 3726 518020 3754
rect 519140 3726 519216 3754
rect 512460 2916 512512 2922
rect 512460 2858 512512 2864
rect 512184 1012 512236 1018
rect 512184 954 512236 960
rect 512472 480 512500 2858
rect 513300 1358 513328 3726
rect 513564 2848 513616 2854
rect 513564 2790 513616 2796
rect 513288 1352 513340 1358
rect 513288 1294 513340 1300
rect 513576 480 513604 2790
rect 514496 1222 514524 3726
rect 515692 2854 515720 3726
rect 516796 2922 516824 3726
rect 516784 2916 516836 2922
rect 516784 2858 516836 2864
rect 515680 2848 515732 2854
rect 515680 2790 515732 2796
rect 517992 1290 518020 3726
rect 515588 1284 515640 1290
rect 515588 1226 515640 1232
rect 517980 1284 518032 1290
rect 517980 1226 518032 1232
rect 514484 1216 514536 1222
rect 514484 1158 514536 1164
rect 514760 1080 514812 1086
rect 514760 1022 514812 1028
rect 514772 480 514800 1022
rect 510038 354 510150 480
rect 509712 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515600 354 515628 1226
rect 517152 1148 517204 1154
rect 517152 1090 517204 1096
rect 517164 480 517192 1090
rect 519188 1086 519216 3726
rect 520200 3726 520272 3754
rect 521440 3754 521468 4012
rect 522636 3754 522664 4012
rect 523740 3754 523768 4012
rect 524936 3754 524964 4012
rect 526040 3754 526068 4012
rect 527236 3754 527264 4012
rect 528432 3754 528460 4012
rect 529536 3754 529564 4012
rect 530732 3754 530760 4012
rect 531836 3754 531864 4012
rect 533032 3754 533060 4012
rect 534228 3754 534256 4012
rect 535332 3754 535360 4012
rect 536528 3754 536556 4012
rect 537632 3754 537660 4012
rect 538828 3754 538856 4012
rect 540024 3754 540052 4012
rect 541128 3754 541156 4012
rect 542324 3754 542352 4012
rect 521440 3726 521516 3754
rect 522636 3726 522712 3754
rect 523740 3726 523816 3754
rect 524936 3726 525012 3754
rect 526040 3726 526116 3754
rect 527236 3726 527312 3754
rect 528432 3726 528508 3754
rect 529536 3726 529612 3754
rect 530732 3726 530808 3754
rect 531836 3726 531912 3754
rect 533032 3726 533108 3754
rect 534228 3726 534304 3754
rect 535332 3726 535408 3754
rect 536528 3726 536604 3754
rect 537632 3726 537708 3754
rect 538828 3726 538904 3754
rect 540024 3726 540100 3754
rect 541128 3726 541204 3754
rect 519544 1352 519596 1358
rect 519544 1294 519596 1300
rect 519176 1080 519228 1086
rect 519176 1022 519228 1028
rect 517980 1012 518032 1018
rect 517980 954 518032 960
rect 515926 354 516038 480
rect 515600 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517992 354 518020 954
rect 519556 480 519584 1294
rect 520200 950 520228 3726
rect 521488 1222 521516 3726
rect 521844 2848 521896 2854
rect 521844 2790 521896 2796
rect 520372 1216 520424 1222
rect 520372 1158 520424 1164
rect 521476 1216 521528 1222
rect 521476 1158 521528 1164
rect 520188 944 520240 950
rect 520188 886 520240 892
rect 518318 354 518430 480
rect 517992 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520384 354 520412 1158
rect 521856 480 521884 2790
rect 522684 1154 522712 3726
rect 523040 2916 523092 2922
rect 523040 2858 523092 2864
rect 522672 1148 522724 1154
rect 522672 1090 522724 1096
rect 523052 480 523080 2858
rect 523788 1018 523816 3726
rect 524984 2922 525012 3726
rect 524972 2916 525024 2922
rect 524972 2858 525024 2864
rect 526088 1358 526116 3726
rect 526076 1352 526128 1358
rect 526076 1294 526128 1300
rect 527284 1290 527312 3726
rect 523868 1284 523920 1290
rect 523868 1226 523920 1232
rect 527272 1284 527324 1290
rect 527272 1226 527324 1232
rect 523776 1012 523828 1018
rect 523776 954 523828 960
rect 520710 354 520822 480
rect 520384 326 520822 354
rect 520710 -960 520822 326
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 523880 354 523908 1226
rect 528480 1222 528508 3726
rect 527824 1216 527876 1222
rect 527824 1158 527876 1164
rect 528468 1216 528520 1222
rect 528468 1158 528520 1164
rect 525432 1080 525484 1086
rect 525432 1022 525484 1028
rect 525444 480 525472 1022
rect 526260 944 526312 950
rect 526260 886 526312 892
rect 524206 354 524318 480
rect 523880 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526272 354 526300 886
rect 527836 480 527864 1158
rect 528652 1148 528704 1154
rect 528652 1090 528704 1096
rect 526598 354 526710 480
rect 526272 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528664 354 528692 1090
rect 529584 950 529612 3726
rect 530780 1154 530808 3726
rect 531320 2916 531372 2922
rect 531320 2858 531372 2864
rect 530768 1148 530820 1154
rect 530768 1090 530820 1096
rect 529940 1012 529992 1018
rect 529940 954 529992 960
rect 529572 944 529624 950
rect 529572 886 529624 892
rect 528990 354 529102 480
rect 528664 326 529102 354
rect 529952 354 529980 954
rect 531332 480 531360 2858
rect 531884 1086 531912 3726
rect 532148 1352 532200 1358
rect 532148 1294 532200 1300
rect 531872 1080 531924 1086
rect 531872 1022 531924 1028
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532160 354 532188 1294
rect 533080 1018 533108 3726
rect 534276 1358 534304 3726
rect 535380 2990 535408 3726
rect 535368 2984 535420 2990
rect 535368 2926 535420 2932
rect 536576 2922 536604 3726
rect 536564 2916 536616 2922
rect 536564 2858 536616 2864
rect 534264 1352 534316 1358
rect 534264 1294 534316 1300
rect 537680 1290 537708 3726
rect 533712 1284 533764 1290
rect 533712 1226 533764 1232
rect 537668 1284 537720 1290
rect 537668 1226 537720 1232
rect 533068 1012 533120 1018
rect 533068 954 533120 960
rect 533724 480 533752 1226
rect 534540 1216 534592 1222
rect 534540 1158 534592 1164
rect 532486 354 532598 480
rect 532160 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534552 354 534580 1158
rect 537208 1148 537260 1154
rect 537208 1090 537260 1096
rect 536104 944 536156 950
rect 536104 886 536156 892
rect 536116 480 536144 886
rect 537220 480 537248 1090
rect 538876 1086 538904 3726
rect 538220 1080 538272 1086
rect 538220 1022 538272 1028
rect 538864 1080 538916 1086
rect 538864 1022 538916 1028
rect 534878 354 534990 480
rect 534552 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 1022
rect 540072 1018 540100 3726
rect 541176 1358 541204 3726
rect 542280 3726 542352 3754
rect 543428 3754 543456 4012
rect 544624 3754 544652 4012
rect 545820 3754 545848 4012
rect 546924 3754 546952 4012
rect 548120 3754 548148 4012
rect 549316 3754 549344 4012
rect 550420 3754 550448 4012
rect 551616 3754 551644 4012
rect 552720 3754 552748 4012
rect 553916 3754 553944 4012
rect 555112 3754 555140 4012
rect 556216 3754 556244 4012
rect 557412 3754 557440 4012
rect 558516 3754 558544 4012
rect 559712 3754 559740 4012
rect 543428 3726 543504 3754
rect 544624 3726 544700 3754
rect 545820 3726 545896 3754
rect 546924 3726 547000 3754
rect 548120 3726 548196 3754
rect 549316 3726 549392 3754
rect 550420 3726 550496 3754
rect 551616 3726 551692 3754
rect 552720 3726 552796 3754
rect 553916 3726 553992 3754
rect 555112 3726 555188 3754
rect 556216 3726 556292 3754
rect 557412 3726 557488 3754
rect 558516 3726 558592 3754
rect 541992 2984 542044 2990
rect 541992 2926 542044 2932
rect 540428 1352 540480 1358
rect 540428 1294 540480 1300
rect 541164 1352 541216 1358
rect 541164 1294 541216 1300
rect 539600 1012 539652 1018
rect 539600 954 539652 960
rect 540060 1012 540112 1018
rect 540060 954 540112 960
rect 539612 480 539640 954
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540440 354 540468 1294
rect 542004 480 542032 2926
rect 542280 1222 542308 3726
rect 543188 2916 543240 2922
rect 543188 2858 543240 2864
rect 542268 1216 542320 1222
rect 542268 1158 542320 1164
rect 543200 480 543228 2858
rect 543476 1154 543504 3726
rect 544672 2922 544700 3726
rect 544660 2916 544712 2922
rect 544660 2858 544712 2864
rect 545868 2854 545896 3726
rect 545856 2848 545908 2854
rect 545856 2790 545908 2796
rect 544384 1284 544436 1290
rect 544384 1226 544436 1232
rect 543464 1148 543516 1154
rect 543464 1090 543516 1096
rect 544396 480 544424 1226
rect 546972 1086 547000 3726
rect 548168 1358 548196 3726
rect 547880 1352 547932 1358
rect 547880 1294 547932 1300
rect 548156 1352 548208 1358
rect 548156 1294 548208 1300
rect 545488 1080 545540 1086
rect 545488 1022 545540 1028
rect 546960 1080 547012 1086
rect 546960 1022 547012 1028
rect 545500 480 545528 1022
rect 546500 1012 546552 1018
rect 546500 954 546552 960
rect 540766 354 540878 480
rect 540440 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 954
rect 547892 480 547920 1294
rect 549364 1290 549392 3726
rect 549352 1284 549404 1290
rect 549352 1226 549404 1232
rect 548708 1216 548760 1222
rect 548708 1158 548760 1164
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548720 354 548748 1158
rect 550468 1154 550496 3726
rect 551468 2916 551520 2922
rect 551468 2858 551520 2864
rect 550272 1148 550324 1154
rect 550272 1090 550324 1096
rect 550456 1148 550508 1154
rect 550456 1090 550508 1096
rect 550284 480 550312 1090
rect 551480 480 551508 2858
rect 551664 1018 551692 3726
rect 552664 2848 552716 2854
rect 552664 2790 552716 2796
rect 551652 1012 551704 1018
rect 551652 954 551704 960
rect 552676 480 552704 2790
rect 552768 882 552796 3726
rect 553964 2922 553992 3726
rect 553952 2916 554004 2922
rect 553952 2858 554004 2864
rect 555160 1358 555188 3726
rect 554780 1352 554832 1358
rect 554780 1294 554832 1300
rect 555148 1352 555200 1358
rect 555148 1294 555200 1300
rect 553768 1080 553820 1086
rect 553768 1022 553820 1028
rect 552756 876 552808 882
rect 552756 818 552808 824
rect 553780 480 553808 1022
rect 549046 354 549158 480
rect 548720 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 1294
rect 556160 1284 556212 1290
rect 556160 1226 556212 1232
rect 556172 480 556200 1226
rect 556264 1222 556292 3726
rect 556252 1216 556304 1222
rect 556252 1158 556304 1164
rect 556988 1148 557040 1154
rect 556988 1090 557040 1096
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 557000 354 557028 1090
rect 557460 626 557488 3726
rect 558564 1154 558592 3726
rect 559668 3726 559740 3754
rect 560908 3754 560936 4012
rect 562012 3754 562040 4012
rect 560908 3726 560984 3754
rect 558552 1148 558604 1154
rect 558552 1090 558604 1096
rect 558552 1012 558604 1018
rect 558552 954 558604 960
rect 557460 610 557580 626
rect 557460 604 557592 610
rect 557460 598 557540 604
rect 557540 546 557592 552
rect 558564 480 558592 954
rect 559668 950 559696 3726
rect 560852 2916 560904 2922
rect 560852 2858 560904 2864
rect 559656 944 559708 950
rect 559656 886 559708 892
rect 559748 876 559800 882
rect 559748 818 559800 824
rect 559760 480 559788 818
rect 560864 480 560892 2858
rect 560956 1086 560984 3726
rect 561968 3726 562040 3754
rect 563208 3754 563236 4012
rect 564312 3754 564340 4012
rect 565508 3754 565536 4012
rect 563208 3726 563284 3754
rect 560944 1080 560996 1086
rect 560944 1022 560996 1028
rect 561968 1018 561996 3726
rect 562048 1352 562100 1358
rect 562048 1294 562100 1300
rect 561956 1012 562008 1018
rect 561956 954 562008 960
rect 562060 480 562088 1294
rect 563256 1290 563284 3726
rect 564268 3726 564340 3754
rect 565464 3726 565536 3754
rect 566704 3754 566732 4012
rect 567808 3754 567836 4012
rect 569004 3754 569032 4012
rect 570108 3754 570136 4012
rect 571304 3754 571332 4012
rect 566704 3726 566780 3754
rect 567808 3726 567884 3754
rect 569004 3726 569080 3754
rect 570108 3726 570184 3754
rect 563244 1284 563296 1290
rect 563244 1226 563296 1232
rect 563152 1216 563204 1222
rect 563152 1158 563204 1164
rect 563164 626 563192 1158
rect 563164 598 563284 626
rect 563256 480 563284 598
rect 557326 354 557438 480
rect 557000 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564268 66 564296 3726
rect 565268 1148 565320 1154
rect 565268 1090 565320 1096
rect 564440 604 564492 610
rect 564440 546 564492 552
rect 564452 480 564480 546
rect 564256 60 564308 66
rect 564256 2 564308 8
rect 564410 -960 564522 480
rect 565280 354 565308 1090
rect 565464 474 565492 3726
rect 566752 1358 566780 3726
rect 566740 1352 566792 1358
rect 566740 1294 566792 1300
rect 567856 1154 567884 3726
rect 569052 1222 569080 3726
rect 569040 1216 569092 1222
rect 569040 1158 569092 1164
rect 567844 1148 567896 1154
rect 567844 1090 567896 1096
rect 567660 1080 567712 1086
rect 567660 1022 567712 1028
rect 566832 944 566884 950
rect 566832 886 566884 892
rect 566844 480 566872 886
rect 565452 468 565504 474
rect 565452 410 565504 416
rect 565606 354 565718 480
rect 565280 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567672 354 567700 1022
rect 570156 1018 570184 3726
rect 571260 3726 571332 3754
rect 572500 3754 572528 4012
rect 573604 3754 573632 4012
rect 574800 3754 574828 4012
rect 575918 3998 576164 4026
rect 572500 3726 572576 3754
rect 573604 3726 573680 3754
rect 574800 3726 574876 3754
rect 570328 1284 570380 1290
rect 570328 1226 570380 1232
rect 568764 1012 568816 1018
rect 568764 954 568816 960
rect 570144 1012 570196 1018
rect 570144 954 570196 960
rect 567998 354 568110 480
rect 567672 326 568110 354
rect 568776 354 568804 954
rect 570340 480 570368 1226
rect 571260 1086 571288 3726
rect 572548 1358 572576 3726
rect 573652 2990 573680 3726
rect 573640 2984 573692 2990
rect 573640 2926 573692 2932
rect 574848 2922 574876 3726
rect 574836 2916 574888 2922
rect 574836 2858 574888 2864
rect 572536 1352 572588 1358
rect 572536 1294 572588 1300
rect 576136 1290 576164 3998
rect 581000 2984 581052 2990
rect 581000 2926 581052 2932
rect 579436 1352 579488 1358
rect 579436 1294 579488 1300
rect 573548 1284 573600 1290
rect 573548 1226 573600 1232
rect 576124 1284 576176 1290
rect 576124 1226 576176 1232
rect 571248 1080 571300 1086
rect 571248 1022 571300 1028
rect 569102 354 569214 480
rect 568776 326 569214 354
rect 567998 -960 568110 326
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571494 82 571606 480
rect 571352 66 571606 82
rect 571340 60 571606 66
rect 571392 54 571606 60
rect 571340 2 571392 8
rect 571494 -960 571606 54
rect 572690 354 572802 480
rect 572904 468 572956 474
rect 572904 410 572956 416
rect 572916 354 572944 410
rect 572690 326 572944 354
rect 573560 354 573588 1226
rect 575940 1216 575992 1222
rect 575940 1158 575992 1164
rect 575112 1148 575164 1154
rect 575112 1090 575164 1096
rect 575124 480 575152 1090
rect 573886 354 573998 480
rect 573560 326 573998 354
rect 572690 -960 572802 326
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 575952 354 575980 1158
rect 578608 1080 578660 1086
rect 578608 1022 578660 1028
rect 577044 1012 577096 1018
rect 577044 954 577096 960
rect 576278 354 576390 480
rect 575952 326 576390 354
rect 577056 354 577084 954
rect 578620 480 578648 1022
rect 577382 354 577494 480
rect 577056 326 577494 354
rect 576278 -960 576390 326
rect 577382 -960 577494 326
rect 578578 -960 578690 480
rect 579448 354 579476 1294
rect 581012 480 581040 2926
rect 582196 2916 582248 2922
rect 582196 2858 582248 2864
rect 582208 480 582236 2858
rect 583392 1284 583444 1290
rect 583392 1226 583444 1232
rect 583404 480 583432 1226
rect 579774 354 579886 480
rect 579448 326 579886 354
rect 579774 -960 579886 326
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 18 698128 74 698184
rect 18 684528 74 684584
rect 579986 683848 580042 683904
rect 578422 682216 578478 682272
rect 2778 680992 2834 681048
rect 2778 671200 2834 671256
rect 579526 670656 579582 670712
rect 579526 666440 579582 666496
rect 3422 664004 3478 664060
rect 3422 658144 3478 658200
rect 578882 650664 578938 650720
rect 18 646992 74 647048
rect 578882 644000 578938 644056
rect 579526 634888 579582 634944
rect 18 632576 74 632632
rect 579618 630808 579674 630864
rect 2778 630264 2834 630320
rect 2778 619112 2834 619168
rect 579526 619112 579582 619168
rect 579618 617480 579674 617536
rect 3422 613252 3478 613308
rect 3422 606056 3478 606112
rect 578882 603336 578938 603392
rect 18 596264 74 596320
rect 578882 590960 578938 591016
rect 578882 587560 578938 587616
rect 18 580488 74 580544
rect 18 579400 74 579456
rect 578882 577632 578938 577688
rect 578882 571784 578938 571840
rect 18 567160 74 567216
rect 578882 564304 578938 564360
rect 2778 562536 2834 562592
rect 578882 556008 578938 556064
rect 2778 553832 2834 553888
rect 18 545536 74 545592
rect 578974 540232 579030 540288
rect 578882 537784 578938 537840
rect 110 528536 166 528592
rect 18 528128 74 528184
rect 578882 524592 578938 524648
rect 110 515344 166 515400
rect 2778 511808 2834 511864
rect 578974 524456 579030 524512
rect 578882 511264 578938 511320
rect 578882 508680 578938 508736
rect 2778 501744 2834 501800
rect 18 494808 74 494864
rect 578974 492768 579030 492824
rect 578882 484608 578938 484664
rect 110 477808 166 477864
rect 18 476040 74 476096
rect 579066 477264 579122 477320
rect 578974 471416 579030 471472
rect 110 463120 166 463176
rect 578882 461488 578938 461544
rect 18 460944 74 461000
rect 18 449792 74 449848
rect 18 444080 74 444136
rect 579066 458088 579122 458144
rect 578974 445576 579030 445632
rect 578882 431568 578938 431624
rect 110 427080 166 427136
rect 570 423580 572 423600
rect 572 423580 624 423600
rect 624 423580 626 423600
rect 570 423544 626 423580
rect 579066 429800 579122 429856
rect 578974 418240 579030 418296
rect 578882 414160 578938 414216
rect 110 411032 166 411088
rect 294 410080 350 410136
rect 578238 398384 578294 398440
rect 294 397976 350 398032
rect 18 393352 74 393408
rect 579066 404912 579122 404968
rect 578974 382472 579030 382528
rect 578882 378392 578938 378448
rect 110 376352 166 376408
rect 18 371864 74 371920
rect 18 359352 74 359408
rect 578882 366832 578938 366888
rect 110 358672 166 358728
rect 578330 351076 578386 351112
rect 578330 351056 578332 351076
rect 578332 351056 578384 351076
rect 578384 351056 578386 351076
rect 18 345888 74 345944
rect 18 342488 74 342544
rect 110 325624 166 325680
rect 18 319776 74 319832
rect 18 308624 74 308680
rect 580262 365064 580318 365120
rect 578974 351872 579030 351928
rect 578974 335416 579030 335472
rect 578882 325216 578938 325272
rect 578882 319504 578938 319560
rect 110 306448 166 306504
rect 578514 303748 578570 303784
rect 578514 303728 578516 303748
rect 578516 303728 578568 303748
rect 578568 303728 578570 303748
rect 18 293664 74 293720
rect 18 291760 74 291816
rect 110 274760 166 274816
rect 18 267416 74 267472
rect 580262 312024 580318 312080
rect 578974 298696 579030 298752
rect 578974 287952 579030 288008
rect 202 257896 258 257952
rect 110 254632 166 254688
rect 578606 256400 578662 256456
rect 579066 272176 579122 272232
rect 578974 245520 579030 245576
rect 202 241440 258 241496
rect 18 240760 74 240816
rect 578882 240624 578938 240680
rect 110 224032 166 224088
rect 18 215192 74 215248
rect 578330 209208 578386 209264
rect 202 207168 258 207224
rect 110 202408 166 202464
rect 18 190168 74 190224
rect 580814 272176 580870 272232
rect 580262 258848 580318 258904
rect 579066 232328 579122 232384
rect 578974 224984 579030 225040
rect 578882 205672 578938 205728
rect 578882 193296 578938 193352
rect 202 189080 258 189136
rect 110 173304 166 173360
rect 18 163376 74 163432
rect 580262 219000 580318 219056
rect 578974 192480 579030 192536
rect 580262 179152 580318 179208
rect 578974 177520 579030 177576
rect 578882 165824 578938 165880
rect 578882 161880 578938 161936
rect 202 156304 258 156360
rect 110 150320 166 150376
rect 18 139440 74 139496
rect 578974 152632 579030 152688
rect 578974 146104 579030 146160
rect 578882 139304 578938 139360
rect 202 137264 258 137320
rect 578882 130192 578938 130248
rect 110 122440 166 122496
rect 18 111152 74 111208
rect 18 105576 74 105632
rect 578974 125976 579030 126032
rect 578974 114552 579030 114608
rect 578882 112784 578938 112840
rect 578974 99456 579030 99512
rect 578882 98776 578938 98832
rect 110 97824 166 97880
rect 110 88712 166 88768
rect 18 85176 74 85232
rect 578882 86128 578938 86184
rect 578882 83000 578938 83056
rect 578882 72936 578938 72992
rect 110 71848 166 71904
rect 294 71304 350 71360
rect 578238 67224 578294 67280
rect 580814 59608 580870 59664
rect 294 59064 350 59120
rect 2778 54848 2834 54904
rect 579526 51448 579582 51504
rect 579526 46280 579582 46336
rect 2778 45464 2834 45520
rect 2042 37848 2098 37904
rect 579526 35672 579582 35728
rect 579618 33088 579674 33144
rect 2042 32408 2098 32464
rect 1306 20984 1362 21040
rect 1306 19352 1362 19408
rect 579618 6568 579674 6624
rect 2778 6432 2834 6488
rect 2778 4120 2834 4176
rect 579526 4120 579582 4176
<< metal3 >>
rect 13 698186 79 698189
rect 13 698184 4110 698186
rect 13 698128 18 698184
rect 74 698128 4110 698184
rect 13 698126 4110 698128
rect 13 698123 79 698126
rect 4050 697948 4110 698126
rect 575920 697918 576410 697978
rect 576350 697914 576410 697918
rect 576350 697854 583586 697914
rect -960 697220 480 697460
rect 583526 697370 583586 697854
rect 583342 697324 583586 697370
rect 583342 697310 584960 697324
rect 583342 697234 583402 697310
rect 583520 697234 584960 697310
rect 583342 697174 584960 697234
rect 583520 697084 584960 697174
rect 13 684586 79 684589
rect 13 684584 122 684586
rect 13 684528 18 684584
rect 74 684528 122 684584
rect 13 684523 122 684528
rect 62 684450 122 684523
rect 62 684404 674 684450
rect -960 684390 674 684404
rect -960 684314 480 684390
rect 614 684314 674 684390
rect -960 684254 674 684314
rect -960 684164 480 684254
rect 579981 683906 580047 683909
rect 583520 683906 584960 683996
rect 579981 683904 584960 683906
rect 579981 683848 579986 683904
rect 580042 683848 584960 683904
rect 579981 683846 584960 683848
rect 579981 683843 580047 683846
rect 583520 683756 584960 683846
rect 578417 682274 578483 682277
rect 576350 682272 578483 682274
rect 576350 682240 578422 682272
rect 575920 682216 578422 682240
rect 578478 682216 578483 682272
rect 575920 682214 578483 682216
rect 575920 682180 576410 682214
rect 578417 682211 578483 682214
rect 2773 681050 2839 681053
rect 2773 681048 3434 681050
rect 2773 680992 2778 681048
rect 2834 681020 3434 681048
rect 2834 680992 4048 681020
rect 2773 680990 4048 680992
rect 2773 680987 2839 680990
rect 3374 680960 4048 680990
rect -960 671258 480 671348
rect 2773 671258 2839 671261
rect -960 671256 2839 671258
rect -960 671200 2778 671256
rect 2834 671200 2839 671256
rect -960 671198 2839 671200
rect -960 671108 480 671198
rect 2773 671195 2839 671198
rect 579521 670714 579587 670717
rect 583520 670714 584960 670804
rect 579521 670712 584960 670714
rect 579521 670656 579526 670712
rect 579582 670656 584960 670712
rect 579521 670654 584960 670656
rect 579521 670651 579587 670654
rect 583520 670564 584960 670654
rect 575920 666498 576410 666502
rect 579521 666498 579587 666501
rect 575920 666496 579587 666498
rect 575920 666442 579526 666496
rect 576350 666440 579526 666442
rect 579582 666440 579587 666496
rect 576350 666438 579587 666440
rect 579521 666435 579587 666438
rect 3417 664062 3483 664065
rect 3417 664060 4048 664062
rect 3417 664004 3422 664060
rect 3478 664004 4048 664060
rect 3417 664002 4048 664004
rect 3417 663999 3483 664002
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect 575920 650722 576410 650764
rect 578877 650722 578943 650725
rect 575920 650720 578943 650722
rect 575920 650704 578882 650720
rect 576350 650664 578882 650704
rect 578938 650664 578943 650720
rect 576350 650662 578943 650664
rect 578877 650659 578943 650662
rect 13 647050 79 647053
rect 3374 647050 4048 647104
rect 13 647048 4048 647050
rect 13 646992 18 647048
rect 74 647044 4048 647048
rect 74 646992 3434 647044
rect 13 646990 3434 646992
rect 13 646987 79 646990
rect -960 644996 480 645236
rect 578877 644058 578943 644061
rect 583520 644058 584960 644148
rect 578877 644056 584960 644058
rect 578877 644000 578882 644056
rect 578938 644000 584960 644056
rect 578877 643998 584960 644000
rect 578877 643995 578943 643998
rect 583520 643908 584960 643998
rect 579521 634946 579587 634949
rect 576350 634944 579587 634946
rect 576350 634904 579526 634944
rect 575920 634888 579526 634904
rect 579582 634888 579587 634944
rect 575920 634886 579587 634888
rect 575920 634844 576410 634886
rect 579521 634883 579587 634886
rect 13 632634 79 632637
rect 13 632632 122 632634
rect 13 632576 18 632632
rect 74 632576 122 632632
rect 13 632571 122 632576
rect 62 632226 122 632571
rect 62 632180 674 632226
rect -960 632166 674 632180
rect -960 632090 480 632166
rect 614 632090 674 632166
rect -960 632030 674 632090
rect -960 631940 480 632030
rect 579613 630866 579679 630869
rect 583520 630866 584960 630956
rect 579613 630864 584960 630866
rect 579613 630808 579618 630864
rect 579674 630808 584960 630864
rect 579613 630806 584960 630808
rect 579613 630803 579679 630806
rect 583520 630716 584960 630806
rect 2773 630322 2839 630325
rect 2773 630320 3434 630322
rect 2773 630264 2778 630320
rect 2834 630268 3434 630320
rect 2834 630264 4048 630268
rect 2773 630262 4048 630264
rect 2773 630259 2839 630262
rect 3374 630208 4048 630262
rect -960 619170 480 619260
rect 2773 619170 2839 619173
rect 579521 619170 579587 619173
rect -960 619168 2839 619170
rect -960 619112 2778 619168
rect 2834 619112 2839 619168
rect 576350 619168 579587 619170
rect 576350 619166 579526 619168
rect -960 619110 2839 619112
rect -960 619020 480 619110
rect 2773 619107 2839 619110
rect 575920 619112 579526 619166
rect 579582 619112 579587 619168
rect 575920 619110 579587 619112
rect 575920 619106 576410 619110
rect 579521 619107 579587 619110
rect 579613 617538 579679 617541
rect 583520 617538 584960 617628
rect 579613 617536 584960 617538
rect 579613 617480 579618 617536
rect 579674 617480 584960 617536
rect 579613 617478 584960 617480
rect 579613 617475 579679 617478
rect 583520 617388 584960 617478
rect 3417 613310 3483 613313
rect 3417 613308 4048 613310
rect 3417 613252 3422 613308
rect 3478 613252 4048 613308
rect 3417 613250 4048 613252
rect 3417 613247 3483 613250
rect -960 606114 480 606204
rect 3417 606114 3483 606117
rect -960 606112 3483 606114
rect -960 606056 3422 606112
rect 3478 606056 3483 606112
rect -960 606054 3483 606056
rect -960 605964 480 606054
rect 3417 606051 3483 606054
rect 583520 604060 584960 604300
rect 575920 603394 576410 603428
rect 578877 603394 578943 603397
rect 575920 603392 578943 603394
rect 575920 603368 578882 603392
rect 576350 603336 578882 603368
rect 578938 603336 578943 603392
rect 576350 603334 578943 603336
rect 578877 603331 578943 603334
rect 13 596322 79 596325
rect 3374 596322 4048 596352
rect 13 596320 4048 596322
rect 13 596264 18 596320
rect 74 596292 4048 596320
rect 74 596264 3434 596292
rect 13 596262 3434 596264
rect 13 596259 79 596262
rect -960 592908 480 593148
rect 578877 591018 578943 591021
rect 583520 591018 584960 591108
rect 578877 591016 584960 591018
rect 578877 590960 578882 591016
rect 578938 590960 584960 591016
rect 578877 590958 584960 590960
rect 578877 590955 578943 590958
rect 583520 590868 584960 590958
rect 575920 587630 576410 587690
rect 576350 587618 576410 587630
rect 578877 587618 578943 587621
rect 576350 587616 578943 587618
rect 576350 587560 578882 587616
rect 578938 587560 578943 587616
rect 576350 587558 578943 587560
rect 578877 587555 578943 587558
rect 13 580546 79 580549
rect 13 580544 122 580546
rect 13 580488 18 580544
rect 74 580488 122 580544
rect 13 580483 122 580488
rect 62 580138 122 580483
rect 62 580092 674 580138
rect -960 580078 674 580092
rect -960 580002 480 580078
rect 614 580002 674 580078
rect -960 579942 674 580002
rect -960 579852 480 579942
rect 13 579458 79 579461
rect 3374 579458 4048 579516
rect 13 579456 4048 579458
rect 13 579400 18 579456
rect 74 579400 3434 579456
rect 13 579398 3434 579400
rect 13 579395 79 579398
rect 578877 577690 578943 577693
rect 583520 577690 584960 577780
rect 578877 577688 584960 577690
rect 578877 577632 578882 577688
rect 578938 577632 584960 577688
rect 578877 577630 584960 577632
rect 578877 577627 578943 577630
rect 583520 577540 584960 577630
rect 578877 571842 578943 571845
rect 576350 571840 578943 571842
rect 576350 571830 578882 571840
rect 575920 571784 578882 571830
rect 578938 571784 578943 571840
rect 575920 571782 578943 571784
rect 575920 571770 576410 571782
rect 578877 571779 578943 571782
rect 13 567218 79 567221
rect 13 567216 122 567218
rect 13 567160 18 567216
rect 74 567160 122 567216
rect 13 567155 122 567160
rect 62 567082 122 567155
rect 62 567036 674 567082
rect -960 567022 674 567036
rect -960 566946 480 567022
rect 614 566946 674 567022
rect -960 566886 674 566946
rect -960 566796 480 566886
rect 578877 564362 578943 564365
rect 583520 564362 584960 564452
rect 578877 564360 584960 564362
rect 578877 564304 578882 564360
rect 578938 564304 584960 564360
rect 578877 564302 584960 564304
rect 578877 564299 578943 564302
rect 583520 564212 584960 564302
rect 2773 562594 2839 562597
rect 2773 562592 3434 562594
rect 2773 562536 2778 562592
rect 2834 562558 3434 562592
rect 2834 562536 4048 562558
rect 2773 562534 4048 562536
rect 2773 562531 2839 562534
rect 3374 562498 4048 562534
rect 575920 556066 576410 556092
rect 578877 556066 578943 556069
rect 575920 556064 578943 556066
rect 575920 556032 578882 556064
rect 576350 556008 578882 556032
rect 578938 556008 578943 556064
rect 576350 556006 578943 556008
rect 578877 556003 578943 556006
rect -960 553890 480 553980
rect 2773 553890 2839 553893
rect -960 553888 2839 553890
rect -960 553832 2778 553888
rect 2834 553832 2839 553888
rect -960 553830 2839 553832
rect -960 553740 480 553830
rect 2773 553827 2839 553830
rect 583520 551020 584960 551260
rect 13 545594 79 545597
rect 3374 545594 4048 545600
rect 13 545592 4048 545594
rect 13 545536 18 545592
rect 74 545540 4048 545592
rect 74 545536 3434 545540
rect 13 545534 3434 545536
rect 13 545531 79 545534
rect -960 540684 480 540924
rect 575920 540294 576410 540354
rect 576350 540290 576410 540294
rect 578969 540290 579035 540293
rect 576350 540288 579035 540290
rect 576350 540232 578974 540288
rect 579030 540232 579035 540288
rect 576350 540230 579035 540232
rect 578969 540227 579035 540230
rect 578877 537842 578943 537845
rect 583520 537842 584960 537932
rect 578877 537840 584960 537842
rect 578877 537784 578882 537840
rect 578938 537784 584960 537840
rect 578877 537782 584960 537784
rect 578877 537779 578943 537782
rect 583520 537692 584960 537782
rect 105 528594 171 528597
rect 3374 528594 4048 528642
rect 105 528592 4048 528594
rect 105 528536 110 528592
rect 166 528582 4048 528592
rect 166 528536 3434 528582
rect 105 528534 3434 528536
rect 105 528531 171 528534
rect 13 528186 79 528189
rect 13 528184 122 528186
rect 13 528128 18 528184
rect 74 528128 122 528184
rect 13 528123 122 528128
rect 62 528050 122 528123
rect 62 528004 674 528050
rect -960 527990 674 528004
rect -960 527914 480 527990
rect 614 527914 674 527990
rect -960 527854 674 527914
rect -960 527764 480 527854
rect 578877 524650 578943 524653
rect 576350 524648 578943 524650
rect 576350 524616 578882 524648
rect 575920 524592 578882 524616
rect 578938 524592 578943 524648
rect 575920 524590 578943 524592
rect 575920 524556 576410 524590
rect 578877 524587 578943 524590
rect 578969 524514 579035 524517
rect 583520 524514 584960 524604
rect 578969 524512 584960 524514
rect 578969 524456 578974 524512
rect 579030 524456 584960 524512
rect 578969 524454 584960 524456
rect 578969 524451 579035 524454
rect 583520 524364 584960 524454
rect 105 515402 171 515405
rect 105 515400 306 515402
rect 105 515344 110 515400
rect 166 515344 306 515400
rect 105 515342 306 515344
rect 105 515339 171 515342
rect 246 514994 306 515342
rect 246 514948 674 514994
rect -960 514934 674 514948
rect -960 514858 480 514934
rect 614 514858 674 514934
rect -960 514798 674 514858
rect -960 514708 480 514798
rect 2773 511866 2839 511869
rect 2773 511864 3434 511866
rect 2773 511808 2778 511864
rect 2834 511808 3434 511864
rect 2773 511806 3434 511808
rect 2773 511803 2839 511806
rect 3374 511746 4048 511806
rect 578877 511322 578943 511325
rect 583520 511322 584960 511412
rect 578877 511320 584960 511322
rect 578877 511264 578882 511320
rect 578938 511264 584960 511320
rect 578877 511262 584960 511264
rect 578877 511259 578943 511262
rect 583520 511172 584960 511262
rect 575920 508738 576410 508756
rect 578877 508738 578943 508741
rect 575920 508736 578943 508738
rect 575920 508696 578882 508736
rect 576350 508680 578882 508696
rect 578938 508680 578943 508736
rect 576350 508678 578943 508680
rect 578877 508675 578943 508678
rect -960 501802 480 501892
rect 2773 501802 2839 501805
rect -960 501800 2839 501802
rect -960 501744 2778 501800
rect 2834 501744 2839 501800
rect -960 501742 2839 501744
rect -960 501652 480 501742
rect 2773 501739 2839 501742
rect 583520 497844 584960 498084
rect 13 494866 79 494869
rect 13 494864 3434 494866
rect 13 494808 18 494864
rect 74 494848 3434 494864
rect 74 494808 4048 494848
rect 13 494806 4048 494808
rect 13 494803 79 494806
rect 3374 494788 4048 494806
rect 575920 492962 576410 493018
rect 575920 492958 576870 492962
rect 576350 492902 576870 492958
rect 576810 492826 576870 492902
rect 578969 492826 579035 492829
rect 576810 492824 579035 492826
rect 576810 492768 578974 492824
rect 579030 492768 579035 492824
rect 576810 492766 579035 492768
rect 578969 492763 579035 492766
rect -960 488596 480 488836
rect 578877 484666 578943 484669
rect 583520 484666 584960 484756
rect 578877 484664 584960 484666
rect 578877 484608 578882 484664
rect 578938 484608 584960 484664
rect 578877 484606 584960 484608
rect 578877 484603 578943 484606
rect 583520 484516 584960 484606
rect 105 477866 171 477869
rect 3374 477866 4048 477890
rect 105 477864 4048 477866
rect 105 477808 110 477864
rect 166 477830 4048 477864
rect 166 477808 3434 477830
rect 105 477806 3434 477808
rect 105 477803 171 477806
rect 579061 477322 579127 477325
rect 576350 477320 579127 477322
rect 576350 477280 579066 477320
rect 575920 477264 579066 477280
rect 579122 477264 579127 477320
rect 575920 477262 579127 477264
rect 575920 477220 576410 477262
rect 579061 477259 579127 477262
rect 13 476098 79 476101
rect 13 476096 122 476098
rect 13 476040 18 476096
rect 74 476040 122 476096
rect 13 476035 122 476040
rect 62 475826 122 476035
rect 62 475780 674 475826
rect -960 475766 674 475780
rect -960 475690 480 475766
rect 614 475690 674 475766
rect -960 475630 674 475690
rect -960 475540 480 475630
rect 578969 471474 579035 471477
rect 583520 471474 584960 471564
rect 578969 471472 584960 471474
rect 578969 471416 578974 471472
rect 579030 471416 584960 471472
rect 578969 471414 584960 471416
rect 578969 471411 579035 471414
rect 583520 471324 584960 471414
rect 105 463178 171 463181
rect 105 463176 306 463178
rect 105 463120 110 463176
rect 166 463120 306 463176
rect 105 463118 306 463120
rect 105 463115 171 463118
rect 246 462770 306 463118
rect 246 462724 674 462770
rect -960 462710 674 462724
rect -960 462634 480 462710
rect 614 462634 674 462710
rect -960 462574 674 462634
rect -960 462484 480 462574
rect 578877 461546 578943 461549
rect 576350 461544 578943 461546
rect 576350 461542 578882 461544
rect 575920 461488 578882 461542
rect 578938 461488 578943 461544
rect 575920 461486 578943 461488
rect 575920 461482 576410 461486
rect 578877 461483 578943 461486
rect 13 461002 79 461005
rect 3374 461002 4048 461054
rect 13 461000 4048 461002
rect 13 460944 18 461000
rect 74 460994 4048 461000
rect 74 460944 3434 460994
rect 13 460942 3434 460944
rect 13 460939 79 460942
rect 579061 458146 579127 458149
rect 583520 458146 584960 458236
rect 579061 458144 584960 458146
rect 579061 458088 579066 458144
rect 579122 458088 584960 458144
rect 579061 458086 584960 458088
rect 579061 458083 579127 458086
rect 583520 457996 584960 458086
rect 13 449850 79 449853
rect 13 449848 122 449850
rect 13 449792 18 449848
rect 74 449792 122 449848
rect 13 449787 122 449792
rect 62 449714 122 449787
rect 62 449668 674 449714
rect -960 449654 674 449668
rect -960 449578 480 449654
rect 614 449578 674 449654
rect -960 449518 674 449578
rect -960 449428 480 449518
rect 575920 445634 576410 445682
rect 578969 445634 579035 445637
rect 575920 445632 579035 445634
rect 575920 445622 578974 445632
rect 576350 445576 578974 445622
rect 579030 445576 579035 445632
rect 576350 445574 579035 445576
rect 578969 445571 579035 445574
rect 583520 444668 584960 444908
rect 13 444138 79 444141
rect 13 444136 3434 444138
rect 13 444080 18 444136
rect 74 444096 3434 444136
rect 74 444080 4048 444096
rect 13 444078 4048 444080
rect 13 444075 79 444078
rect 3374 444036 4048 444078
rect -960 436508 480 436748
rect 578877 431626 578943 431629
rect 583520 431626 584960 431716
rect 578877 431624 584960 431626
rect 578877 431568 578882 431624
rect 578938 431568 584960 431624
rect 578877 431566 584960 431568
rect 578877 431563 578943 431566
rect 583520 431476 584960 431566
rect 575920 429884 576410 429944
rect 576350 429858 576410 429884
rect 579061 429858 579127 429861
rect 576350 429856 579127 429858
rect 576350 429800 579066 429856
rect 579122 429800 579127 429856
rect 576350 429798 579127 429800
rect 579061 429795 579127 429798
rect 105 427138 171 427141
rect 105 427136 4048 427138
rect 105 427080 110 427136
rect 166 427080 4048 427136
rect 105 427078 4048 427080
rect 105 427075 171 427078
rect -960 423602 480 423692
rect 565 423602 631 423605
rect -960 423600 631 423602
rect -960 423544 570 423600
rect 626 423544 631 423600
rect -960 423542 631 423544
rect -960 423452 480 423542
rect 565 423539 631 423542
rect 578969 418298 579035 418301
rect 583520 418298 584960 418388
rect 578969 418296 584960 418298
rect 578969 418240 578974 418296
rect 579030 418240 584960 418296
rect 578969 418238 584960 418240
rect 578969 418235 579035 418238
rect 583520 418148 584960 418238
rect 578877 414218 578943 414221
rect 576350 414216 578943 414218
rect 576350 414206 578882 414216
rect 575920 414160 578882 414206
rect 578938 414160 578943 414216
rect 575920 414158 578943 414160
rect 575920 414146 576410 414158
rect 578877 414155 578943 414158
rect 105 411090 171 411093
rect 105 411088 306 411090
rect 105 411032 110 411088
rect 166 411032 306 411088
rect 105 411030 306 411032
rect 105 411027 171 411030
rect 246 410682 306 411030
rect 246 410636 674 410682
rect -960 410622 674 410636
rect -960 410546 480 410622
rect 614 410546 674 410622
rect -960 410486 674 410546
rect -960 410396 480 410486
rect 289 410138 355 410141
rect 3374 410138 4048 410180
rect 289 410136 4048 410138
rect 289 410080 294 410136
rect 350 410120 4048 410136
rect 350 410080 3434 410120
rect 289 410078 3434 410080
rect 289 410075 355 410078
rect 579061 404970 579127 404973
rect 583520 404970 584960 405060
rect 579061 404968 584960 404970
rect 579061 404912 579066 404968
rect 579122 404912 584960 404968
rect 579061 404910 584960 404912
rect 579061 404907 579127 404910
rect 583520 404820 584960 404910
rect 575920 398442 576410 398468
rect 578233 398442 578299 398445
rect 575920 398440 578299 398442
rect 575920 398408 578238 398440
rect 576350 398384 578238 398408
rect 578294 398384 578299 398440
rect 576350 398382 578299 398384
rect 578233 398379 578299 398382
rect 289 398034 355 398037
rect 246 398032 355 398034
rect 246 397976 294 398032
rect 350 397976 355 398032
rect 246 397971 355 397976
rect 246 397626 306 397971
rect 246 397580 674 397626
rect -960 397566 674 397580
rect -960 397490 480 397566
rect 614 397490 674 397566
rect -960 397430 674 397490
rect -960 397340 480 397430
rect 13 393410 79 393413
rect 13 393408 3802 393410
rect 13 393352 18 393408
rect 74 393352 3802 393408
rect 13 393350 3802 393352
rect 13 393347 79 393350
rect 3742 393344 3802 393350
rect 3742 393284 4048 393344
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 575920 382548 576410 382608
rect 576350 382530 576410 382548
rect 578969 382530 579035 382533
rect 576350 382528 579035 382530
rect 576350 382472 578974 382528
rect 579030 382472 579035 382528
rect 576350 382470 579035 382472
rect 578969 382467 579035 382470
rect 578877 378450 578943 378453
rect 583520 378450 584960 378540
rect 578877 378448 584960 378450
rect 578877 378392 578882 378448
rect 578938 378392 584960 378448
rect 578877 378390 584960 378392
rect 578877 378387 578943 378390
rect 583520 378300 584960 378390
rect 105 376410 171 376413
rect 105 376408 3434 376410
rect 105 376352 110 376408
rect 166 376386 3434 376408
rect 166 376352 4048 376386
rect 105 376350 4048 376352
rect 105 376347 171 376350
rect 3374 376326 4048 376350
rect 13 371922 79 371925
rect 13 371920 122 371922
rect 13 371864 18 371920
rect 74 371864 122 371920
rect 13 371859 122 371864
rect 62 371514 122 371859
rect 62 371468 674 371514
rect -960 371454 674 371468
rect -960 371378 480 371454
rect 614 371378 674 371454
rect -960 371318 674 371378
rect -960 371228 480 371318
rect 578877 366890 578943 366893
rect 576350 366888 578943 366890
rect 576350 366870 578882 366888
rect 575920 366832 578882 366870
rect 578938 366832 578943 366888
rect 575920 366830 578943 366832
rect 575920 366810 576410 366830
rect 578877 366827 578943 366830
rect 580257 365122 580323 365125
rect 583520 365122 584960 365212
rect 580257 365120 584960 365122
rect 580257 365064 580262 365120
rect 580318 365064 584960 365120
rect 580257 365062 584960 365064
rect 580257 365059 580323 365062
rect 583520 364972 584960 365062
rect 13 359410 79 359413
rect 3374 359410 4048 359428
rect 13 359408 4048 359410
rect 13 359352 18 359408
rect 74 359368 4048 359408
rect 74 359352 3434 359368
rect 13 359350 3434 359352
rect 13 359347 79 359350
rect 105 358730 171 358733
rect 105 358728 306 358730
rect 105 358672 110 358728
rect 166 358672 306 358728
rect 105 358670 306 358672
rect 105 358667 171 358670
rect 246 358594 306 358670
rect 246 358548 674 358594
rect -960 358534 674 358548
rect -960 358458 480 358534
rect 614 358458 674 358534
rect -960 358398 674 358458
rect -960 358308 480 358398
rect 578969 351930 579035 351933
rect 583520 351930 584960 352020
rect 578969 351928 584960 351930
rect 578969 351872 578974 351928
rect 579030 351872 584960 351928
rect 578969 351870 584960 351872
rect 578969 351867 579035 351870
rect 583520 351780 584960 351870
rect 575920 351114 576410 351132
rect 578325 351114 578391 351117
rect 575920 351112 578391 351114
rect 575920 351072 578330 351112
rect 576350 351056 578330 351072
rect 578386 351056 578391 351112
rect 576350 351054 578391 351056
rect 578325 351051 578391 351054
rect 13 345946 79 345949
rect 13 345944 122 345946
rect 13 345888 18 345944
rect 74 345888 122 345944
rect 13 345883 122 345888
rect 62 345538 122 345883
rect 62 345492 674 345538
rect -960 345478 674 345492
rect -960 345402 480 345478
rect 614 345402 674 345478
rect -960 345342 674 345402
rect -960 345252 480 345342
rect 13 342546 79 342549
rect 3374 342546 4048 342592
rect 13 342544 4048 342546
rect 13 342488 18 342544
rect 74 342532 4048 342544
rect 74 342488 3434 342532
rect 13 342486 3434 342488
rect 13 342483 79 342486
rect 583520 338452 584960 338692
rect 578969 335474 579035 335477
rect 576350 335472 579035 335474
rect 576350 335416 578974 335472
rect 579030 335416 579035 335472
rect 576350 335414 579035 335416
rect 576350 335394 576410 335414
rect 578969 335411 579035 335414
rect 575920 335334 576410 335394
rect -960 332196 480 332436
rect 105 325682 171 325685
rect 105 325680 3434 325682
rect 105 325624 110 325680
rect 166 325634 3434 325680
rect 166 325624 4048 325634
rect 105 325622 4048 325624
rect 105 325619 171 325622
rect 3374 325574 4048 325622
rect 578877 325274 578943 325277
rect 583520 325274 584960 325364
rect 578877 325272 584960 325274
rect 578877 325216 578882 325272
rect 578938 325216 584960 325272
rect 578877 325214 584960 325216
rect 578877 325211 578943 325214
rect 583520 325124 584960 325214
rect 13 319834 79 319837
rect 13 319832 122 319834
rect 13 319776 18 319832
rect 74 319776 122 319832
rect 13 319771 122 319776
rect 62 319426 122 319771
rect 578877 319562 578943 319565
rect 576350 319560 578943 319562
rect 576350 319534 578882 319560
rect 575920 319504 578882 319534
rect 578938 319504 578943 319560
rect 575920 319502 578943 319504
rect 575920 319474 576410 319502
rect 578877 319499 578943 319502
rect 62 319380 674 319426
rect -960 319366 674 319380
rect -960 319290 480 319366
rect 614 319290 674 319366
rect -960 319230 674 319290
rect -960 319140 480 319230
rect 580257 312082 580323 312085
rect 583520 312082 584960 312172
rect 580257 312080 584960 312082
rect 580257 312024 580262 312080
rect 580318 312024 584960 312080
rect 580257 312022 584960 312024
rect 580257 312019 580323 312022
rect 583520 311932 584960 312022
rect 13 308682 79 308685
rect 13 308680 3434 308682
rect 13 308624 18 308680
rect 74 308676 3434 308680
rect 74 308624 4048 308676
rect 13 308622 4048 308624
rect 13 308619 79 308622
rect 3374 308616 4048 308622
rect 105 306506 171 306509
rect 62 306504 171 306506
rect 62 306448 110 306504
rect 166 306448 171 306504
rect 62 306443 171 306448
rect 62 306370 122 306443
rect 62 306324 674 306370
rect -960 306310 674 306324
rect -960 306234 480 306310
rect 614 306234 674 306310
rect -960 306174 674 306234
rect -960 306084 480 306174
rect 575920 303786 576410 303796
rect 578509 303786 578575 303789
rect 575920 303784 578575 303786
rect 575920 303736 578514 303784
rect 576350 303728 578514 303736
rect 578570 303728 578575 303784
rect 576350 303726 578575 303728
rect 578509 303723 578575 303726
rect 578969 298754 579035 298757
rect 583520 298754 584960 298844
rect 578969 298752 584960 298754
rect 578969 298696 578974 298752
rect 579030 298696 584960 298752
rect 578969 298694 584960 298696
rect 578969 298691 579035 298694
rect 583520 298604 584960 298694
rect 13 293722 79 293725
rect 13 293720 122 293722
rect 13 293664 18 293720
rect 74 293664 122 293720
rect 13 293659 122 293664
rect 62 293314 122 293659
rect 62 293268 674 293314
rect -960 293254 674 293268
rect -960 293178 480 293254
rect 614 293178 674 293254
rect -960 293118 674 293178
rect -960 293028 480 293118
rect 13 291818 79 291821
rect 3374 291818 4048 291840
rect 13 291816 4048 291818
rect 13 291760 18 291816
rect 74 291780 4048 291816
rect 74 291760 3434 291780
rect 13 291758 3434 291760
rect 13 291755 79 291758
rect 575920 288010 576410 288058
rect 578969 288010 579035 288013
rect 575920 288008 579035 288010
rect 575920 287998 578974 288008
rect 576350 287952 578974 287998
rect 579030 287952 579035 288008
rect 576350 287950 579035 287952
rect 578969 287947 579035 287950
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 3742 274822 4048 274882
rect 105 274818 171 274821
rect 3742 274818 3802 274822
rect 105 274816 3802 274818
rect 105 274760 110 274816
rect 166 274760 3802 274816
rect 105 274758 3802 274760
rect 105 274755 171 274758
rect 575920 272260 576410 272320
rect 576350 272234 576410 272260
rect 579061 272234 579127 272237
rect 576350 272232 579127 272234
rect 576350 272176 579066 272232
rect 579122 272176 579127 272232
rect 576350 272174 579127 272176
rect 579061 272171 579127 272174
rect 580809 272234 580875 272237
rect 583520 272234 584960 272324
rect 580809 272232 584960 272234
rect 580809 272176 580814 272232
rect 580870 272176 584960 272232
rect 580809 272174 584960 272176
rect 580809 272171 580875 272174
rect 583520 272084 584960 272174
rect 13 267474 79 267477
rect 13 267472 122 267474
rect 13 267416 18 267472
rect 74 267416 122 267472
rect 13 267411 122 267416
rect 62 267338 122 267411
rect 62 267292 674 267338
rect -960 267278 674 267292
rect -960 267202 480 267278
rect 614 267202 674 267278
rect -960 267142 674 267202
rect -960 267052 480 267142
rect 580257 258906 580323 258909
rect 583520 258906 584960 258996
rect 580257 258904 584960 258906
rect 580257 258848 580262 258904
rect 580318 258848 584960 258904
rect 580257 258846 584960 258848
rect 580257 258843 580323 258846
rect 583520 258756 584960 258846
rect 197 257954 263 257957
rect 197 257952 3434 257954
rect 197 257896 202 257952
rect 258 257924 3434 257952
rect 258 257896 4048 257924
rect 197 257894 4048 257896
rect 197 257891 263 257894
rect 3374 257864 4048 257894
rect 575920 256458 576410 256460
rect 578601 256458 578667 256461
rect 575920 256456 578667 256458
rect 575920 256400 578606 256456
rect 578662 256400 578667 256456
rect 576350 256398 578667 256400
rect 578601 256395 578667 256398
rect 105 254690 171 254693
rect 105 254688 306 254690
rect 105 254632 110 254688
rect 166 254632 306 254688
rect 105 254630 306 254632
rect 105 254627 171 254630
rect 246 254282 306 254630
rect 246 254236 674 254282
rect -960 254222 674 254236
rect -960 254146 480 254222
rect 614 254146 674 254222
rect -960 254086 674 254146
rect -960 253996 480 254086
rect 578969 245578 579035 245581
rect 583520 245578 584960 245668
rect 578969 245576 584960 245578
rect 578969 245520 578974 245576
rect 579030 245520 584960 245576
rect 578969 245518 584960 245520
rect 578969 245515 579035 245518
rect 583520 245428 584960 245518
rect 197 241498 263 241501
rect 197 241496 306 241498
rect 197 241440 202 241496
rect 258 241440 306 241496
rect 197 241435 306 241440
rect 246 241226 306 241435
rect 246 241180 674 241226
rect -960 241166 674 241180
rect -960 241090 480 241166
rect 614 241090 674 241166
rect -960 241030 674 241090
rect -960 240940 480 241030
rect 3374 240906 4048 240966
rect 13 240818 79 240821
rect 3374 240818 3434 240906
rect 13 240816 3434 240818
rect 13 240760 18 240816
rect 74 240760 3434 240816
rect 13 240758 3434 240760
rect 13 240755 79 240758
rect 575920 240682 576410 240722
rect 578877 240682 578943 240685
rect 575920 240680 578943 240682
rect 575920 240662 578882 240680
rect 576350 240624 578882 240662
rect 578938 240624 578943 240680
rect 576350 240622 578943 240624
rect 578877 240619 578943 240622
rect 579061 232386 579127 232389
rect 583520 232386 584960 232476
rect 579061 232384 584960 232386
rect 579061 232328 579066 232384
rect 579122 232328 584960 232384
rect 579061 232326 584960 232328
rect 579061 232323 579127 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 578969 225042 579035 225045
rect 576350 225040 579035 225042
rect 576350 224984 578974 225040
rect 579030 224984 579035 225040
rect 575920 224982 579035 224984
rect 575920 224924 576410 224982
rect 578969 224979 579035 224982
rect 105 224090 171 224093
rect 3374 224090 4048 224130
rect 105 224088 4048 224090
rect 105 224032 110 224088
rect 166 224070 4048 224088
rect 166 224032 3434 224070
rect 105 224030 3434 224032
rect 105 224027 171 224030
rect 580257 219058 580323 219061
rect 583520 219058 584960 219148
rect 580257 219056 584960 219058
rect 580257 219000 580262 219056
rect 580318 219000 584960 219056
rect 580257 218998 584960 219000
rect 580257 218995 580323 218998
rect 583520 218908 584960 218998
rect 13 215250 79 215253
rect 13 215248 122 215250
rect 13 215192 18 215248
rect 74 215192 122 215248
rect 13 215187 122 215192
rect 62 215114 122 215187
rect 62 215068 674 215114
rect -960 215054 674 215068
rect -960 214978 480 215054
rect 614 214978 674 215054
rect -960 214918 674 214978
rect -960 214828 480 214918
rect 578325 209266 578391 209269
rect 576350 209264 578391 209266
rect 576350 209246 578330 209264
rect 575920 209208 578330 209246
rect 578386 209208 578391 209264
rect 575920 209206 578391 209208
rect 575920 209186 576410 209206
rect 578325 209203 578391 209206
rect 197 207226 263 207229
rect 197 207224 3434 207226
rect 197 207168 202 207224
rect 258 207172 3434 207224
rect 258 207168 4048 207172
rect 197 207166 4048 207168
rect 197 207163 263 207166
rect 3374 207112 4048 207166
rect 578877 205730 578943 205733
rect 583520 205730 584960 205820
rect 578877 205728 584960 205730
rect 578877 205672 578882 205728
rect 578938 205672 584960 205728
rect 578877 205670 584960 205672
rect 578877 205667 578943 205670
rect 583520 205580 584960 205670
rect 105 202466 171 202469
rect 105 202464 306 202466
rect 105 202408 110 202464
rect 166 202408 306 202464
rect 105 202406 306 202408
rect 105 202403 171 202406
rect 246 202058 306 202406
rect 246 202012 674 202058
rect -960 201998 674 202012
rect -960 201922 480 201998
rect 614 201922 674 201998
rect -960 201862 674 201922
rect -960 201772 480 201862
rect 575920 193354 576410 193386
rect 578877 193354 578943 193357
rect 575920 193352 578943 193354
rect 575920 193326 578882 193352
rect 576350 193296 578882 193326
rect 578938 193296 578943 193352
rect 576350 193294 578943 193296
rect 578877 193291 578943 193294
rect 578969 192538 579035 192541
rect 583520 192538 584960 192628
rect 578969 192536 584960 192538
rect 578969 192480 578974 192536
rect 579030 192480 584960 192536
rect 578969 192478 584960 192480
rect 578969 192475 579035 192478
rect 583520 192388 584960 192478
rect 13 190226 79 190229
rect 13 190224 3434 190226
rect 13 190168 18 190224
rect 74 190214 3434 190224
rect 74 190168 4048 190214
rect 13 190166 4048 190168
rect 13 190163 79 190166
rect 3374 190154 4048 190166
rect 197 189138 263 189141
rect 197 189136 306 189138
rect 197 189080 202 189136
rect 258 189080 306 189136
rect 197 189075 306 189080
rect 246 189002 306 189075
rect 246 188956 674 189002
rect -960 188942 674 188956
rect -960 188866 480 188942
rect 614 188866 674 188942
rect -960 188806 674 188866
rect -960 188716 480 188806
rect 580257 179210 580323 179213
rect 583520 179210 584960 179300
rect 580257 179208 584960 179210
rect 580257 179152 580262 179208
rect 580318 179152 584960 179208
rect 580257 179150 584960 179152
rect 580257 179147 580323 179150
rect 583520 179060 584960 179150
rect 575920 177588 576410 177648
rect 576350 177578 576410 177588
rect 578969 177578 579035 177581
rect 576350 177576 579035 177578
rect 576350 177520 578974 177576
rect 579030 177520 579035 177576
rect 576350 177518 579035 177520
rect 578969 177515 579035 177518
rect -960 175796 480 176036
rect 105 173362 171 173365
rect 3374 173362 4048 173378
rect 105 173360 4048 173362
rect 105 173304 110 173360
rect 166 173318 4048 173360
rect 166 173304 3434 173318
rect 105 173302 3434 173304
rect 105 173299 171 173302
rect 578877 165882 578943 165885
rect 583520 165882 584960 165972
rect 578877 165880 584960 165882
rect 578877 165824 578882 165880
rect 578938 165824 584960 165880
rect 578877 165822 584960 165824
rect 578877 165819 578943 165822
rect 583520 165732 584960 165822
rect 13 163434 79 163437
rect 13 163432 122 163434
rect 13 163376 18 163432
rect 74 163376 122 163432
rect 13 163371 122 163376
rect 62 163026 122 163371
rect 62 162980 674 163026
rect -960 162966 674 162980
rect -960 162890 480 162966
rect 614 162890 674 162966
rect -960 162830 674 162890
rect -960 162740 480 162830
rect 578877 161938 578943 161941
rect 576350 161936 578943 161938
rect 576350 161910 578882 161936
rect 575920 161880 578882 161910
rect 578938 161880 578943 161936
rect 575920 161878 578943 161880
rect 575920 161850 576410 161878
rect 578877 161875 578943 161878
rect 197 156362 263 156365
rect 3374 156362 4048 156420
rect 197 156360 4048 156362
rect 197 156304 202 156360
rect 258 156304 3434 156360
rect 197 156302 3434 156304
rect 197 156299 263 156302
rect 578969 152690 579035 152693
rect 583520 152690 584960 152780
rect 578969 152688 584960 152690
rect 578969 152632 578974 152688
rect 579030 152632 584960 152688
rect 578969 152630 584960 152632
rect 578969 152627 579035 152630
rect 583520 152540 584960 152630
rect 105 150378 171 150381
rect 105 150376 306 150378
rect 105 150320 110 150376
rect 166 150320 306 150376
rect 105 150318 306 150320
rect 105 150315 171 150318
rect 246 149970 306 150318
rect 246 149924 674 149970
rect -960 149910 674 149924
rect -960 149834 480 149910
rect 614 149834 674 149910
rect -960 149774 674 149834
rect -960 149684 480 149774
rect 575920 146162 576410 146172
rect 578969 146162 579035 146165
rect 575920 146160 579035 146162
rect 575920 146112 578974 146160
rect 576350 146104 578974 146112
rect 579030 146104 579035 146160
rect 576350 146102 579035 146104
rect 578969 146099 579035 146102
rect 13 139498 79 139501
rect 13 139496 3434 139498
rect 13 139440 18 139496
rect 74 139462 3434 139496
rect 74 139440 4048 139462
rect 13 139438 4048 139440
rect 13 139435 79 139438
rect 3374 139402 4048 139438
rect 578877 139362 578943 139365
rect 583520 139362 584960 139452
rect 578877 139360 584960 139362
rect 578877 139304 578882 139360
rect 578938 139304 584960 139360
rect 578877 139302 584960 139304
rect 578877 139299 578943 139302
rect 583520 139212 584960 139302
rect 197 137322 263 137325
rect 197 137320 306 137322
rect 197 137264 202 137320
rect 258 137264 306 137320
rect 197 137259 306 137264
rect 246 136914 306 137259
rect 246 136868 674 136914
rect -960 136854 674 136868
rect -960 136778 480 136854
rect 614 136778 674 136854
rect -960 136718 674 136778
rect -960 136628 480 136718
rect 575920 130252 576410 130312
rect 576350 130250 576410 130252
rect 578877 130250 578943 130253
rect 576350 130248 578943 130250
rect 576350 130192 578882 130248
rect 578938 130192 578943 130248
rect 576350 130190 578943 130192
rect 578877 130187 578943 130190
rect 578969 126034 579035 126037
rect 583520 126034 584960 126124
rect 578969 126032 584960 126034
rect 578969 125976 578974 126032
rect 579030 125976 584960 126032
rect 578969 125974 584960 125976
rect 578969 125971 579035 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 105 122498 171 122501
rect 3374 122498 4048 122504
rect 105 122496 4048 122498
rect 105 122440 110 122496
rect 166 122444 4048 122496
rect 166 122440 3434 122444
rect 105 122438 3434 122440
rect 105 122435 171 122438
rect 578969 114610 579035 114613
rect 576350 114608 579035 114610
rect 576350 114574 578974 114608
rect 575920 114552 578974 114574
rect 579030 114552 579035 114608
rect 575920 114550 579035 114552
rect 575920 114514 576410 114550
rect 578969 114547 579035 114550
rect 578877 112842 578943 112845
rect 583520 112842 584960 112932
rect 578877 112840 584960 112842
rect 578877 112784 578882 112840
rect 578938 112784 584960 112840
rect 578877 112782 584960 112784
rect 578877 112779 578943 112782
rect 583520 112692 584960 112782
rect 13 111210 79 111213
rect 13 111208 122 111210
rect 13 111152 18 111208
rect 74 111152 122 111208
rect 13 111147 122 111152
rect 62 110802 122 111147
rect 62 110756 674 110802
rect -960 110742 674 110756
rect -960 110666 480 110742
rect 614 110666 674 110742
rect -960 110606 674 110666
rect -960 110516 480 110606
rect 13 105634 79 105637
rect 3374 105634 4048 105668
rect 13 105632 4048 105634
rect 13 105576 18 105632
rect 74 105608 4048 105632
rect 74 105576 3434 105608
rect 13 105574 3434 105576
rect 13 105571 79 105574
rect 578969 99514 579035 99517
rect 583520 99514 584960 99604
rect 578969 99512 584960 99514
rect 578969 99456 578974 99512
rect 579030 99456 584960 99512
rect 578969 99454 584960 99456
rect 578969 99451 579035 99454
rect 583520 99364 584960 99454
rect 575920 98834 576410 98836
rect 578877 98834 578943 98837
rect 575920 98832 578943 98834
rect 575920 98776 578882 98832
rect 578938 98776 578943 98832
rect 576350 98774 578943 98776
rect 578877 98771 578943 98774
rect 105 97882 171 97885
rect 105 97880 306 97882
rect 105 97824 110 97880
rect 166 97824 306 97880
rect 105 97822 306 97824
rect 105 97819 171 97822
rect 246 97746 306 97822
rect 246 97700 674 97746
rect -960 97686 674 97700
rect -960 97610 480 97686
rect 614 97610 674 97686
rect -960 97550 674 97610
rect -960 97460 480 97550
rect 105 88770 171 88773
rect 105 88768 3434 88770
rect 105 88712 110 88768
rect 166 88712 3434 88768
rect 105 88710 3434 88712
rect 105 88707 171 88710
rect 3374 88650 4048 88710
rect 578877 86186 578943 86189
rect 583520 86186 584960 86276
rect 578877 86184 584960 86186
rect 578877 86128 578882 86184
rect 578938 86128 584960 86184
rect 578877 86126 584960 86128
rect 578877 86123 578943 86126
rect 583520 86036 584960 86126
rect 13 85234 79 85237
rect 13 85232 122 85234
rect 13 85176 18 85232
rect 74 85176 122 85232
rect 13 85171 122 85176
rect 62 84826 122 85171
rect 62 84780 674 84826
rect -960 84766 674 84780
rect -960 84690 480 84766
rect 614 84690 674 84766
rect -960 84630 674 84690
rect -960 84540 480 84630
rect 575920 83058 576410 83098
rect 578877 83058 578943 83061
rect 575920 83056 578943 83058
rect 575920 83038 578882 83056
rect 576350 83000 578882 83038
rect 578938 83000 578943 83056
rect 576350 82998 578943 83000
rect 578877 82995 578943 82998
rect 578877 72994 578943 72997
rect 583520 72994 584960 73084
rect 578877 72992 584960 72994
rect 578877 72936 578882 72992
rect 578938 72936 584960 72992
rect 578877 72934 584960 72936
rect 578877 72931 578943 72934
rect 583520 72844 584960 72934
rect 105 71906 171 71909
rect 62 71904 171 71906
rect 62 71848 110 71904
rect 166 71848 171 71904
rect 62 71843 171 71848
rect 62 71770 122 71843
rect 62 71724 674 71770
rect -960 71710 674 71724
rect -960 71634 480 71710
rect 614 71634 674 71710
rect -960 71574 674 71634
rect 3374 71692 4048 71752
rect -960 71484 480 71574
rect 289 71362 355 71365
rect 3374 71362 3434 71692
rect 289 71360 3434 71362
rect 289 71304 294 71360
rect 350 71304 3434 71360
rect 289 71302 3434 71304
rect 289 71299 355 71302
rect 578233 67282 578299 67285
rect 576350 67280 578299 67282
rect 576350 67238 578238 67280
rect 575920 67224 578238 67238
rect 578294 67224 578299 67280
rect 575920 67222 578299 67224
rect 575920 67178 576410 67222
rect 578233 67219 578299 67222
rect 580809 59666 580875 59669
rect 583520 59666 584960 59756
rect 580809 59664 584960 59666
rect 580809 59608 580814 59664
rect 580870 59608 584960 59664
rect 580809 59606 584960 59608
rect 580809 59603 580875 59606
rect 583520 59516 584960 59606
rect 289 59122 355 59125
rect 246 59120 355 59122
rect 246 59064 294 59120
rect 350 59064 355 59120
rect 246 59059 355 59064
rect 246 58714 306 59059
rect 246 58668 674 58714
rect -960 58654 674 58668
rect -960 58578 480 58654
rect 614 58578 674 58654
rect -960 58518 674 58578
rect -960 58428 480 58518
rect 2773 54906 2839 54909
rect 3374 54906 4048 54916
rect 2773 54904 4048 54906
rect 2773 54848 2778 54904
rect 2834 54856 4048 54904
rect 2834 54848 3434 54856
rect 2773 54846 3434 54848
rect 2773 54843 2839 54846
rect 579521 51506 579587 51509
rect 576350 51504 579587 51506
rect 576350 51500 579526 51504
rect 575920 51448 579526 51500
rect 579582 51448 579587 51504
rect 575920 51446 579587 51448
rect 575920 51440 576410 51446
rect 579521 51443 579587 51446
rect 579521 46338 579587 46341
rect 583520 46338 584960 46428
rect 579521 46336 584960 46338
rect 579521 46280 579526 46336
rect 579582 46280 584960 46336
rect 579521 46278 584960 46280
rect 579521 46275 579587 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 2773 45522 2839 45525
rect -960 45520 2839 45522
rect -960 45464 2778 45520
rect 2834 45464 2839 45520
rect -960 45462 2839 45464
rect -960 45372 480 45462
rect 2773 45459 2839 45462
rect 2037 37906 2103 37909
rect 3374 37906 4048 37958
rect 2037 37904 4048 37906
rect 2037 37848 2042 37904
rect 2098 37898 4048 37904
rect 2098 37848 3434 37898
rect 2037 37846 3434 37848
rect 2037 37843 2103 37846
rect 575920 35730 576410 35762
rect 579521 35730 579587 35733
rect 575920 35728 579587 35730
rect 575920 35702 579526 35728
rect 576350 35672 579526 35702
rect 579582 35672 579587 35728
rect 576350 35670 579587 35672
rect 579521 35667 579587 35670
rect 579613 33146 579679 33149
rect 583520 33146 584960 33236
rect 579613 33144 584960 33146
rect 579613 33088 579618 33144
rect 579674 33088 584960 33144
rect 579613 33086 584960 33088
rect 579613 33083 579679 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2037 32466 2103 32469
rect -960 32464 2103 32466
rect -960 32408 2042 32464
rect 2098 32408 2103 32464
rect -960 32406 2103 32408
rect -960 32316 480 32406
rect 2037 32403 2103 32406
rect 1301 21042 1367 21045
rect 1301 21040 3434 21042
rect 1301 20984 1306 21040
rect 1362 21000 3434 21040
rect 1362 20984 4048 21000
rect 1301 20982 4048 20984
rect 1301 20979 1367 20982
rect 3374 20940 4048 20982
rect 575920 19964 576410 20024
rect 576350 19954 576410 19964
rect 576350 19894 576870 19954
rect 576810 19818 576870 19894
rect 583520 19818 584960 19908
rect 576810 19758 584960 19818
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 1301 19410 1367 19413
rect -960 19408 1367 19410
rect -960 19352 1306 19408
rect 1362 19352 1367 19408
rect -960 19350 1367 19352
rect -960 19260 480 19350
rect 1301 19347 1367 19350
rect 579613 6626 579679 6629
rect 583520 6626 584960 6716
rect 579613 6624 584960 6626
rect -960 6490 480 6580
rect 579613 6568 579618 6624
rect 579674 6568 584960 6624
rect 579613 6566 584960 6568
rect 579613 6563 579679 6566
rect 2773 6490 2839 6493
rect -960 6488 2839 6490
rect -960 6432 2778 6488
rect 2834 6432 2839 6488
rect 583520 6476 584960 6566
rect -960 6430 2839 6432
rect -960 6340 480 6430
rect 2773 6427 2839 6430
rect 2773 4178 2839 4181
rect 579521 4178 579587 4181
rect 2773 4176 3802 4178
rect 2773 4120 2778 4176
rect 2834 4164 3802 4176
rect 576166 4176 579587 4178
rect 576166 4164 579526 4176
rect 2834 4120 4048 4164
rect 2773 4118 4048 4120
rect 2773 4115 2839 4118
rect 3742 4104 4048 4118
rect 575920 4120 579526 4164
rect 579582 4120 579587 4176
rect 575920 4118 579587 4120
rect 575920 4104 576226 4118
rect 579521 4115 579587 4118
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 700008 2414 704282
rect 5514 700008 6134 706202
rect 9234 700008 9854 708122
rect 12954 700008 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 700008 20414 705242
rect 23514 700008 24134 707162
rect 27234 700008 27854 709082
rect 30954 700008 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 700008 38414 704282
rect 41514 700008 42134 706202
rect 45234 700008 45854 708122
rect 48954 700008 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 700008 56414 705242
rect 59514 700008 60134 707162
rect 63234 700008 63854 709082
rect 66954 700008 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 700008 74414 704282
rect 77514 700008 78134 706202
rect 81234 700008 81854 708122
rect 84954 700008 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 700008 92414 705242
rect 95514 700008 96134 707162
rect 99234 700008 99854 709082
rect 102954 700008 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 700008 110414 704282
rect 113514 700008 114134 706202
rect 117234 700008 117854 708122
rect 120954 700008 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 700008 128414 705242
rect 131514 700008 132134 707162
rect 135234 700008 135854 709082
rect 138954 700008 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 700008 146414 704282
rect 149514 700008 150134 706202
rect 153234 700008 153854 708122
rect 156954 700008 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 700008 164414 705242
rect 167514 700008 168134 707162
rect 171234 700008 171854 709082
rect 174954 700008 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 700008 182414 704282
rect 185514 700008 186134 706202
rect 189234 700008 189854 708122
rect 192954 700008 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 700008 200414 705242
rect 203514 700008 204134 707162
rect 207234 700008 207854 709082
rect 210954 700008 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 700008 218414 704282
rect 221514 700008 222134 706202
rect 225234 700008 225854 708122
rect 228954 700008 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 700008 236414 705242
rect 239514 700008 240134 707162
rect 243234 700008 243854 709082
rect 246954 700008 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 700008 254414 704282
rect 257514 700008 258134 706202
rect 261234 700008 261854 708122
rect 264954 700008 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 700008 272414 705242
rect 275514 700008 276134 707162
rect 279234 700008 279854 709082
rect 282954 700008 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 700008 290414 704282
rect 293514 700008 294134 706202
rect 297234 700008 297854 708122
rect 300954 700008 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 700008 308414 705242
rect 311514 700008 312134 707162
rect 315234 700008 315854 709082
rect 318954 700008 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 700008 326414 704282
rect 329514 700008 330134 706202
rect 333234 700008 333854 708122
rect 336954 700008 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 700008 344414 705242
rect 347514 700008 348134 707162
rect 351234 700008 351854 709082
rect 354954 700008 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 700008 362414 704282
rect 365514 700008 366134 706202
rect 369234 700008 369854 708122
rect 372954 700008 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 700008 380414 705242
rect 383514 700008 384134 707162
rect 387234 700008 387854 709082
rect 390954 700008 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 700008 398414 704282
rect 401514 700008 402134 706202
rect 405234 700008 405854 708122
rect 408954 700008 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 700008 416414 705242
rect 419514 700008 420134 707162
rect 423234 700008 423854 709082
rect 426954 700008 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 700008 434414 704282
rect 437514 700008 438134 706202
rect 441234 700008 441854 708122
rect 444954 700008 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 700008 452414 705242
rect 455514 700008 456134 707162
rect 459234 700008 459854 709082
rect 462954 700008 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 700008 470414 704282
rect 473514 700008 474134 706202
rect 477234 700008 477854 708122
rect 480954 700008 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 700008 488414 705242
rect 491514 700008 492134 707162
rect 495234 700008 495854 709082
rect 498954 700008 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 700008 506414 704282
rect 509514 700008 510134 706202
rect 513234 700008 513854 708122
rect 516954 700008 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 700008 524414 705242
rect 527514 700008 528134 707162
rect 531234 700008 531854 709082
rect 534954 700008 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 700008 542414 704282
rect 545514 700008 546134 706202
rect 549234 700008 549854 708122
rect 552954 700008 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 700008 560414 705242
rect 563514 700008 564134 707162
rect 567234 700008 567854 709082
rect 570954 700008 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 700008 578414 704282
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect 9084 687454 9704 687486
rect 9084 687218 9116 687454
rect 9352 687218 9436 687454
rect 9672 687218 9704 687454
rect 9084 687134 9704 687218
rect 9084 686898 9116 687134
rect 9352 686898 9436 687134
rect 9672 686898 9704 687134
rect 9084 686866 9704 686898
rect 31200 687454 31872 687486
rect 31200 687218 31258 687454
rect 31494 687218 31578 687454
rect 31814 687218 31872 687454
rect 31200 687134 31872 687218
rect 31200 686898 31258 687134
rect 31494 686898 31578 687134
rect 31814 686898 31872 687134
rect 31200 686866 31872 686898
rect 58400 687454 59072 687486
rect 58400 687218 58458 687454
rect 58694 687218 58778 687454
rect 59014 687218 59072 687454
rect 58400 687134 59072 687218
rect 58400 686898 58458 687134
rect 58694 686898 58778 687134
rect 59014 686898 59072 687134
rect 58400 686866 59072 686898
rect 85600 687454 86272 687486
rect 85600 687218 85658 687454
rect 85894 687218 85978 687454
rect 86214 687218 86272 687454
rect 85600 687134 86272 687218
rect 85600 686898 85658 687134
rect 85894 686898 85978 687134
rect 86214 686898 86272 687134
rect 85600 686866 86272 686898
rect 112800 687454 113472 687486
rect 112800 687218 112858 687454
rect 113094 687218 113178 687454
rect 113414 687218 113472 687454
rect 112800 687134 113472 687218
rect 112800 686898 112858 687134
rect 113094 686898 113178 687134
rect 113414 686898 113472 687134
rect 112800 686866 113472 686898
rect 140000 687454 140672 687486
rect 140000 687218 140058 687454
rect 140294 687218 140378 687454
rect 140614 687218 140672 687454
rect 140000 687134 140672 687218
rect 140000 686898 140058 687134
rect 140294 686898 140378 687134
rect 140614 686898 140672 687134
rect 140000 686866 140672 686898
rect 167200 687454 167872 687486
rect 167200 687218 167258 687454
rect 167494 687218 167578 687454
rect 167814 687218 167872 687454
rect 167200 687134 167872 687218
rect 167200 686898 167258 687134
rect 167494 686898 167578 687134
rect 167814 686898 167872 687134
rect 167200 686866 167872 686898
rect 194400 687454 195072 687486
rect 194400 687218 194458 687454
rect 194694 687218 194778 687454
rect 195014 687218 195072 687454
rect 194400 687134 195072 687218
rect 194400 686898 194458 687134
rect 194694 686898 194778 687134
rect 195014 686898 195072 687134
rect 194400 686866 195072 686898
rect 221600 687454 222272 687486
rect 221600 687218 221658 687454
rect 221894 687218 221978 687454
rect 222214 687218 222272 687454
rect 221600 687134 222272 687218
rect 221600 686898 221658 687134
rect 221894 686898 221978 687134
rect 222214 686898 222272 687134
rect 221600 686866 222272 686898
rect 248800 687454 249472 687486
rect 248800 687218 248858 687454
rect 249094 687218 249178 687454
rect 249414 687218 249472 687454
rect 248800 687134 249472 687218
rect 248800 686898 248858 687134
rect 249094 686898 249178 687134
rect 249414 686898 249472 687134
rect 248800 686866 249472 686898
rect 276000 687454 276672 687486
rect 276000 687218 276058 687454
rect 276294 687218 276378 687454
rect 276614 687218 276672 687454
rect 276000 687134 276672 687218
rect 276000 686898 276058 687134
rect 276294 686898 276378 687134
rect 276614 686898 276672 687134
rect 276000 686866 276672 686898
rect 303200 687454 303872 687486
rect 303200 687218 303258 687454
rect 303494 687218 303578 687454
rect 303814 687218 303872 687454
rect 303200 687134 303872 687218
rect 303200 686898 303258 687134
rect 303494 686898 303578 687134
rect 303814 686898 303872 687134
rect 303200 686866 303872 686898
rect 330400 687454 331072 687486
rect 330400 687218 330458 687454
rect 330694 687218 330778 687454
rect 331014 687218 331072 687454
rect 330400 687134 331072 687218
rect 330400 686898 330458 687134
rect 330694 686898 330778 687134
rect 331014 686898 331072 687134
rect 330400 686866 331072 686898
rect 357600 687454 358272 687486
rect 357600 687218 357658 687454
rect 357894 687218 357978 687454
rect 358214 687218 358272 687454
rect 357600 687134 358272 687218
rect 357600 686898 357658 687134
rect 357894 686898 357978 687134
rect 358214 686898 358272 687134
rect 357600 686866 358272 686898
rect 384800 687454 385472 687486
rect 384800 687218 384858 687454
rect 385094 687218 385178 687454
rect 385414 687218 385472 687454
rect 384800 687134 385472 687218
rect 384800 686898 384858 687134
rect 385094 686898 385178 687134
rect 385414 686898 385472 687134
rect 384800 686866 385472 686898
rect 412000 687454 412672 687486
rect 412000 687218 412058 687454
rect 412294 687218 412378 687454
rect 412614 687218 412672 687454
rect 412000 687134 412672 687218
rect 412000 686898 412058 687134
rect 412294 686898 412378 687134
rect 412614 686898 412672 687134
rect 412000 686866 412672 686898
rect 439200 687454 439872 687486
rect 439200 687218 439258 687454
rect 439494 687218 439578 687454
rect 439814 687218 439872 687454
rect 439200 687134 439872 687218
rect 439200 686898 439258 687134
rect 439494 686898 439578 687134
rect 439814 686898 439872 687134
rect 439200 686866 439872 686898
rect 466400 687454 467072 687486
rect 466400 687218 466458 687454
rect 466694 687218 466778 687454
rect 467014 687218 467072 687454
rect 466400 687134 467072 687218
rect 466400 686898 466458 687134
rect 466694 686898 466778 687134
rect 467014 686898 467072 687134
rect 466400 686866 467072 686898
rect 493600 687454 494272 687486
rect 493600 687218 493658 687454
rect 493894 687218 493978 687454
rect 494214 687218 494272 687454
rect 493600 687134 494272 687218
rect 493600 686898 493658 687134
rect 493894 686898 493978 687134
rect 494214 686898 494272 687134
rect 493600 686866 494272 686898
rect 520800 687454 521472 687486
rect 520800 687218 520858 687454
rect 521094 687218 521178 687454
rect 521414 687218 521472 687454
rect 520800 687134 521472 687218
rect 520800 686898 520858 687134
rect 521094 686898 521178 687134
rect 521414 686898 521472 687134
rect 520800 686866 521472 686898
rect 548000 687454 548672 687486
rect 548000 687218 548058 687454
rect 548294 687218 548378 687454
rect 548614 687218 548672 687454
rect 548000 687134 548672 687218
rect 548000 686898 548058 687134
rect 548294 686898 548378 687134
rect 548614 686898 548672 687134
rect 548000 686866 548672 686898
rect 570260 687454 570880 687486
rect 570260 687218 570292 687454
rect 570528 687218 570612 687454
rect 570848 687218 570880 687454
rect 570260 687134 570880 687218
rect 570260 686898 570292 687134
rect 570528 686898 570612 687134
rect 570848 686898 570880 687134
rect 570260 686866 570880 686898
rect 7844 669454 8464 669486
rect 7844 669218 7876 669454
rect 8112 669218 8196 669454
rect 8432 669218 8464 669454
rect 7844 669134 8464 669218
rect 7844 668898 7876 669134
rect 8112 668898 8196 669134
rect 8432 668898 8464 669134
rect 7844 668866 8464 668898
rect 17600 669454 18272 669486
rect 17600 669218 17658 669454
rect 17894 669218 17978 669454
rect 18214 669218 18272 669454
rect 17600 669134 18272 669218
rect 17600 668898 17658 669134
rect 17894 668898 17978 669134
rect 18214 668898 18272 669134
rect 17600 668866 18272 668898
rect 44800 669454 45472 669486
rect 44800 669218 44858 669454
rect 45094 669218 45178 669454
rect 45414 669218 45472 669454
rect 44800 669134 45472 669218
rect 44800 668898 44858 669134
rect 45094 668898 45178 669134
rect 45414 668898 45472 669134
rect 44800 668866 45472 668898
rect 72000 669454 72672 669486
rect 72000 669218 72058 669454
rect 72294 669218 72378 669454
rect 72614 669218 72672 669454
rect 72000 669134 72672 669218
rect 72000 668898 72058 669134
rect 72294 668898 72378 669134
rect 72614 668898 72672 669134
rect 72000 668866 72672 668898
rect 99200 669454 99872 669486
rect 99200 669218 99258 669454
rect 99494 669218 99578 669454
rect 99814 669218 99872 669454
rect 99200 669134 99872 669218
rect 99200 668898 99258 669134
rect 99494 668898 99578 669134
rect 99814 668898 99872 669134
rect 99200 668866 99872 668898
rect 126400 669454 127072 669486
rect 126400 669218 126458 669454
rect 126694 669218 126778 669454
rect 127014 669218 127072 669454
rect 126400 669134 127072 669218
rect 126400 668898 126458 669134
rect 126694 668898 126778 669134
rect 127014 668898 127072 669134
rect 126400 668866 127072 668898
rect 153600 669454 154272 669486
rect 153600 669218 153658 669454
rect 153894 669218 153978 669454
rect 154214 669218 154272 669454
rect 153600 669134 154272 669218
rect 153600 668898 153658 669134
rect 153894 668898 153978 669134
rect 154214 668898 154272 669134
rect 153600 668866 154272 668898
rect 180800 669454 181472 669486
rect 180800 669218 180858 669454
rect 181094 669218 181178 669454
rect 181414 669218 181472 669454
rect 180800 669134 181472 669218
rect 180800 668898 180858 669134
rect 181094 668898 181178 669134
rect 181414 668898 181472 669134
rect 180800 668866 181472 668898
rect 208000 669454 208672 669486
rect 208000 669218 208058 669454
rect 208294 669218 208378 669454
rect 208614 669218 208672 669454
rect 208000 669134 208672 669218
rect 208000 668898 208058 669134
rect 208294 668898 208378 669134
rect 208614 668898 208672 669134
rect 208000 668866 208672 668898
rect 235200 669454 235872 669486
rect 235200 669218 235258 669454
rect 235494 669218 235578 669454
rect 235814 669218 235872 669454
rect 235200 669134 235872 669218
rect 235200 668898 235258 669134
rect 235494 668898 235578 669134
rect 235814 668898 235872 669134
rect 235200 668866 235872 668898
rect 262400 669454 263072 669486
rect 262400 669218 262458 669454
rect 262694 669218 262778 669454
rect 263014 669218 263072 669454
rect 262400 669134 263072 669218
rect 262400 668898 262458 669134
rect 262694 668898 262778 669134
rect 263014 668898 263072 669134
rect 262400 668866 263072 668898
rect 289600 669454 290272 669486
rect 289600 669218 289658 669454
rect 289894 669218 289978 669454
rect 290214 669218 290272 669454
rect 289600 669134 290272 669218
rect 289600 668898 289658 669134
rect 289894 668898 289978 669134
rect 290214 668898 290272 669134
rect 289600 668866 290272 668898
rect 316800 669454 317472 669486
rect 316800 669218 316858 669454
rect 317094 669218 317178 669454
rect 317414 669218 317472 669454
rect 316800 669134 317472 669218
rect 316800 668898 316858 669134
rect 317094 668898 317178 669134
rect 317414 668898 317472 669134
rect 316800 668866 317472 668898
rect 344000 669454 344672 669486
rect 344000 669218 344058 669454
rect 344294 669218 344378 669454
rect 344614 669218 344672 669454
rect 344000 669134 344672 669218
rect 344000 668898 344058 669134
rect 344294 668898 344378 669134
rect 344614 668898 344672 669134
rect 344000 668866 344672 668898
rect 371200 669454 371872 669486
rect 371200 669218 371258 669454
rect 371494 669218 371578 669454
rect 371814 669218 371872 669454
rect 371200 669134 371872 669218
rect 371200 668898 371258 669134
rect 371494 668898 371578 669134
rect 371814 668898 371872 669134
rect 371200 668866 371872 668898
rect 398400 669454 399072 669486
rect 398400 669218 398458 669454
rect 398694 669218 398778 669454
rect 399014 669218 399072 669454
rect 398400 669134 399072 669218
rect 398400 668898 398458 669134
rect 398694 668898 398778 669134
rect 399014 668898 399072 669134
rect 398400 668866 399072 668898
rect 425600 669454 426272 669486
rect 425600 669218 425658 669454
rect 425894 669218 425978 669454
rect 426214 669218 426272 669454
rect 425600 669134 426272 669218
rect 425600 668898 425658 669134
rect 425894 668898 425978 669134
rect 426214 668898 426272 669134
rect 425600 668866 426272 668898
rect 452800 669454 453472 669486
rect 452800 669218 452858 669454
rect 453094 669218 453178 669454
rect 453414 669218 453472 669454
rect 452800 669134 453472 669218
rect 452800 668898 452858 669134
rect 453094 668898 453178 669134
rect 453414 668898 453472 669134
rect 452800 668866 453472 668898
rect 480000 669454 480672 669486
rect 480000 669218 480058 669454
rect 480294 669218 480378 669454
rect 480614 669218 480672 669454
rect 480000 669134 480672 669218
rect 480000 668898 480058 669134
rect 480294 668898 480378 669134
rect 480614 668898 480672 669134
rect 480000 668866 480672 668898
rect 507200 669454 507872 669486
rect 507200 669218 507258 669454
rect 507494 669218 507578 669454
rect 507814 669218 507872 669454
rect 507200 669134 507872 669218
rect 507200 668898 507258 669134
rect 507494 668898 507578 669134
rect 507814 668898 507872 669134
rect 507200 668866 507872 668898
rect 534400 669454 535072 669486
rect 534400 669218 534458 669454
rect 534694 669218 534778 669454
rect 535014 669218 535072 669454
rect 534400 669134 535072 669218
rect 534400 668898 534458 669134
rect 534694 668898 534778 669134
rect 535014 668898 535072 669134
rect 534400 668866 535072 668898
rect 561600 669454 562272 669486
rect 561600 669218 561658 669454
rect 561894 669218 561978 669454
rect 562214 669218 562272 669454
rect 561600 669134 562272 669218
rect 561600 668898 561658 669134
rect 561894 668898 561978 669134
rect 562214 668898 562272 669134
rect 561600 668866 562272 668898
rect 571500 669454 572120 669486
rect 571500 669218 571532 669454
rect 571768 669218 571852 669454
rect 572088 669218 572120 669454
rect 571500 669134 572120 669218
rect 571500 668898 571532 669134
rect 571768 668898 571852 669134
rect 572088 668898 572120 669134
rect 571500 668866 572120 668898
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect 9084 651454 9704 651486
rect 9084 651218 9116 651454
rect 9352 651218 9436 651454
rect 9672 651218 9704 651454
rect 9084 651134 9704 651218
rect 9084 650898 9116 651134
rect 9352 650898 9436 651134
rect 9672 650898 9704 651134
rect 9084 650866 9704 650898
rect 31200 651454 31872 651486
rect 31200 651218 31258 651454
rect 31494 651218 31578 651454
rect 31814 651218 31872 651454
rect 31200 651134 31872 651218
rect 31200 650898 31258 651134
rect 31494 650898 31578 651134
rect 31814 650898 31872 651134
rect 31200 650866 31872 650898
rect 58400 651454 59072 651486
rect 58400 651218 58458 651454
rect 58694 651218 58778 651454
rect 59014 651218 59072 651454
rect 58400 651134 59072 651218
rect 58400 650898 58458 651134
rect 58694 650898 58778 651134
rect 59014 650898 59072 651134
rect 58400 650866 59072 650898
rect 85600 651454 86272 651486
rect 85600 651218 85658 651454
rect 85894 651218 85978 651454
rect 86214 651218 86272 651454
rect 85600 651134 86272 651218
rect 85600 650898 85658 651134
rect 85894 650898 85978 651134
rect 86214 650898 86272 651134
rect 85600 650866 86272 650898
rect 112800 651454 113472 651486
rect 112800 651218 112858 651454
rect 113094 651218 113178 651454
rect 113414 651218 113472 651454
rect 112800 651134 113472 651218
rect 112800 650898 112858 651134
rect 113094 650898 113178 651134
rect 113414 650898 113472 651134
rect 112800 650866 113472 650898
rect 140000 651454 140672 651486
rect 140000 651218 140058 651454
rect 140294 651218 140378 651454
rect 140614 651218 140672 651454
rect 140000 651134 140672 651218
rect 140000 650898 140058 651134
rect 140294 650898 140378 651134
rect 140614 650898 140672 651134
rect 140000 650866 140672 650898
rect 167200 651454 167872 651486
rect 167200 651218 167258 651454
rect 167494 651218 167578 651454
rect 167814 651218 167872 651454
rect 167200 651134 167872 651218
rect 167200 650898 167258 651134
rect 167494 650898 167578 651134
rect 167814 650898 167872 651134
rect 167200 650866 167872 650898
rect 194400 651454 195072 651486
rect 194400 651218 194458 651454
rect 194694 651218 194778 651454
rect 195014 651218 195072 651454
rect 194400 651134 195072 651218
rect 194400 650898 194458 651134
rect 194694 650898 194778 651134
rect 195014 650898 195072 651134
rect 194400 650866 195072 650898
rect 221600 651454 222272 651486
rect 221600 651218 221658 651454
rect 221894 651218 221978 651454
rect 222214 651218 222272 651454
rect 221600 651134 222272 651218
rect 221600 650898 221658 651134
rect 221894 650898 221978 651134
rect 222214 650898 222272 651134
rect 221600 650866 222272 650898
rect 248800 651454 249472 651486
rect 248800 651218 248858 651454
rect 249094 651218 249178 651454
rect 249414 651218 249472 651454
rect 248800 651134 249472 651218
rect 248800 650898 248858 651134
rect 249094 650898 249178 651134
rect 249414 650898 249472 651134
rect 248800 650866 249472 650898
rect 276000 651454 276672 651486
rect 276000 651218 276058 651454
rect 276294 651218 276378 651454
rect 276614 651218 276672 651454
rect 276000 651134 276672 651218
rect 276000 650898 276058 651134
rect 276294 650898 276378 651134
rect 276614 650898 276672 651134
rect 276000 650866 276672 650898
rect 303200 651454 303872 651486
rect 303200 651218 303258 651454
rect 303494 651218 303578 651454
rect 303814 651218 303872 651454
rect 303200 651134 303872 651218
rect 303200 650898 303258 651134
rect 303494 650898 303578 651134
rect 303814 650898 303872 651134
rect 303200 650866 303872 650898
rect 330400 651454 331072 651486
rect 330400 651218 330458 651454
rect 330694 651218 330778 651454
rect 331014 651218 331072 651454
rect 330400 651134 331072 651218
rect 330400 650898 330458 651134
rect 330694 650898 330778 651134
rect 331014 650898 331072 651134
rect 330400 650866 331072 650898
rect 357600 651454 358272 651486
rect 357600 651218 357658 651454
rect 357894 651218 357978 651454
rect 358214 651218 358272 651454
rect 357600 651134 358272 651218
rect 357600 650898 357658 651134
rect 357894 650898 357978 651134
rect 358214 650898 358272 651134
rect 357600 650866 358272 650898
rect 384800 651454 385472 651486
rect 384800 651218 384858 651454
rect 385094 651218 385178 651454
rect 385414 651218 385472 651454
rect 384800 651134 385472 651218
rect 384800 650898 384858 651134
rect 385094 650898 385178 651134
rect 385414 650898 385472 651134
rect 384800 650866 385472 650898
rect 412000 651454 412672 651486
rect 412000 651218 412058 651454
rect 412294 651218 412378 651454
rect 412614 651218 412672 651454
rect 412000 651134 412672 651218
rect 412000 650898 412058 651134
rect 412294 650898 412378 651134
rect 412614 650898 412672 651134
rect 412000 650866 412672 650898
rect 439200 651454 439872 651486
rect 439200 651218 439258 651454
rect 439494 651218 439578 651454
rect 439814 651218 439872 651454
rect 439200 651134 439872 651218
rect 439200 650898 439258 651134
rect 439494 650898 439578 651134
rect 439814 650898 439872 651134
rect 439200 650866 439872 650898
rect 466400 651454 467072 651486
rect 466400 651218 466458 651454
rect 466694 651218 466778 651454
rect 467014 651218 467072 651454
rect 466400 651134 467072 651218
rect 466400 650898 466458 651134
rect 466694 650898 466778 651134
rect 467014 650898 467072 651134
rect 466400 650866 467072 650898
rect 493600 651454 494272 651486
rect 493600 651218 493658 651454
rect 493894 651218 493978 651454
rect 494214 651218 494272 651454
rect 493600 651134 494272 651218
rect 493600 650898 493658 651134
rect 493894 650898 493978 651134
rect 494214 650898 494272 651134
rect 493600 650866 494272 650898
rect 520800 651454 521472 651486
rect 520800 651218 520858 651454
rect 521094 651218 521178 651454
rect 521414 651218 521472 651454
rect 520800 651134 521472 651218
rect 520800 650898 520858 651134
rect 521094 650898 521178 651134
rect 521414 650898 521472 651134
rect 520800 650866 521472 650898
rect 548000 651454 548672 651486
rect 548000 651218 548058 651454
rect 548294 651218 548378 651454
rect 548614 651218 548672 651454
rect 548000 651134 548672 651218
rect 548000 650898 548058 651134
rect 548294 650898 548378 651134
rect 548614 650898 548672 651134
rect 548000 650866 548672 650898
rect 570260 651454 570880 651486
rect 570260 651218 570292 651454
rect 570528 651218 570612 651454
rect 570848 651218 570880 651454
rect 570260 651134 570880 651218
rect 570260 650898 570292 651134
rect 570528 650898 570612 651134
rect 570848 650898 570880 651134
rect 570260 650866 570880 650898
rect 7844 633454 8464 633486
rect 7844 633218 7876 633454
rect 8112 633218 8196 633454
rect 8432 633218 8464 633454
rect 7844 633134 8464 633218
rect 7844 632898 7876 633134
rect 8112 632898 8196 633134
rect 8432 632898 8464 633134
rect 7844 632866 8464 632898
rect 17600 633454 18272 633486
rect 17600 633218 17658 633454
rect 17894 633218 17978 633454
rect 18214 633218 18272 633454
rect 17600 633134 18272 633218
rect 17600 632898 17658 633134
rect 17894 632898 17978 633134
rect 18214 632898 18272 633134
rect 17600 632866 18272 632898
rect 44800 633454 45472 633486
rect 44800 633218 44858 633454
rect 45094 633218 45178 633454
rect 45414 633218 45472 633454
rect 44800 633134 45472 633218
rect 44800 632898 44858 633134
rect 45094 632898 45178 633134
rect 45414 632898 45472 633134
rect 44800 632866 45472 632898
rect 72000 633454 72672 633486
rect 72000 633218 72058 633454
rect 72294 633218 72378 633454
rect 72614 633218 72672 633454
rect 72000 633134 72672 633218
rect 72000 632898 72058 633134
rect 72294 632898 72378 633134
rect 72614 632898 72672 633134
rect 72000 632866 72672 632898
rect 99200 633454 99872 633486
rect 99200 633218 99258 633454
rect 99494 633218 99578 633454
rect 99814 633218 99872 633454
rect 99200 633134 99872 633218
rect 99200 632898 99258 633134
rect 99494 632898 99578 633134
rect 99814 632898 99872 633134
rect 99200 632866 99872 632898
rect 126400 633454 127072 633486
rect 126400 633218 126458 633454
rect 126694 633218 126778 633454
rect 127014 633218 127072 633454
rect 126400 633134 127072 633218
rect 126400 632898 126458 633134
rect 126694 632898 126778 633134
rect 127014 632898 127072 633134
rect 126400 632866 127072 632898
rect 153600 633454 154272 633486
rect 153600 633218 153658 633454
rect 153894 633218 153978 633454
rect 154214 633218 154272 633454
rect 153600 633134 154272 633218
rect 153600 632898 153658 633134
rect 153894 632898 153978 633134
rect 154214 632898 154272 633134
rect 153600 632866 154272 632898
rect 180800 633454 181472 633486
rect 180800 633218 180858 633454
rect 181094 633218 181178 633454
rect 181414 633218 181472 633454
rect 180800 633134 181472 633218
rect 180800 632898 180858 633134
rect 181094 632898 181178 633134
rect 181414 632898 181472 633134
rect 180800 632866 181472 632898
rect 208000 633454 208672 633486
rect 208000 633218 208058 633454
rect 208294 633218 208378 633454
rect 208614 633218 208672 633454
rect 208000 633134 208672 633218
rect 208000 632898 208058 633134
rect 208294 632898 208378 633134
rect 208614 632898 208672 633134
rect 208000 632866 208672 632898
rect 235200 633454 235872 633486
rect 235200 633218 235258 633454
rect 235494 633218 235578 633454
rect 235814 633218 235872 633454
rect 235200 633134 235872 633218
rect 235200 632898 235258 633134
rect 235494 632898 235578 633134
rect 235814 632898 235872 633134
rect 235200 632866 235872 632898
rect 262400 633454 263072 633486
rect 262400 633218 262458 633454
rect 262694 633218 262778 633454
rect 263014 633218 263072 633454
rect 262400 633134 263072 633218
rect 262400 632898 262458 633134
rect 262694 632898 262778 633134
rect 263014 632898 263072 633134
rect 262400 632866 263072 632898
rect 289600 633454 290272 633486
rect 289600 633218 289658 633454
rect 289894 633218 289978 633454
rect 290214 633218 290272 633454
rect 289600 633134 290272 633218
rect 289600 632898 289658 633134
rect 289894 632898 289978 633134
rect 290214 632898 290272 633134
rect 289600 632866 290272 632898
rect 316800 633454 317472 633486
rect 316800 633218 316858 633454
rect 317094 633218 317178 633454
rect 317414 633218 317472 633454
rect 316800 633134 317472 633218
rect 316800 632898 316858 633134
rect 317094 632898 317178 633134
rect 317414 632898 317472 633134
rect 316800 632866 317472 632898
rect 344000 633454 344672 633486
rect 344000 633218 344058 633454
rect 344294 633218 344378 633454
rect 344614 633218 344672 633454
rect 344000 633134 344672 633218
rect 344000 632898 344058 633134
rect 344294 632898 344378 633134
rect 344614 632898 344672 633134
rect 344000 632866 344672 632898
rect 371200 633454 371872 633486
rect 371200 633218 371258 633454
rect 371494 633218 371578 633454
rect 371814 633218 371872 633454
rect 371200 633134 371872 633218
rect 371200 632898 371258 633134
rect 371494 632898 371578 633134
rect 371814 632898 371872 633134
rect 371200 632866 371872 632898
rect 398400 633454 399072 633486
rect 398400 633218 398458 633454
rect 398694 633218 398778 633454
rect 399014 633218 399072 633454
rect 398400 633134 399072 633218
rect 398400 632898 398458 633134
rect 398694 632898 398778 633134
rect 399014 632898 399072 633134
rect 398400 632866 399072 632898
rect 425600 633454 426272 633486
rect 425600 633218 425658 633454
rect 425894 633218 425978 633454
rect 426214 633218 426272 633454
rect 425600 633134 426272 633218
rect 425600 632898 425658 633134
rect 425894 632898 425978 633134
rect 426214 632898 426272 633134
rect 425600 632866 426272 632898
rect 452800 633454 453472 633486
rect 452800 633218 452858 633454
rect 453094 633218 453178 633454
rect 453414 633218 453472 633454
rect 452800 633134 453472 633218
rect 452800 632898 452858 633134
rect 453094 632898 453178 633134
rect 453414 632898 453472 633134
rect 452800 632866 453472 632898
rect 480000 633454 480672 633486
rect 480000 633218 480058 633454
rect 480294 633218 480378 633454
rect 480614 633218 480672 633454
rect 480000 633134 480672 633218
rect 480000 632898 480058 633134
rect 480294 632898 480378 633134
rect 480614 632898 480672 633134
rect 480000 632866 480672 632898
rect 507200 633454 507872 633486
rect 507200 633218 507258 633454
rect 507494 633218 507578 633454
rect 507814 633218 507872 633454
rect 507200 633134 507872 633218
rect 507200 632898 507258 633134
rect 507494 632898 507578 633134
rect 507814 632898 507872 633134
rect 507200 632866 507872 632898
rect 534400 633454 535072 633486
rect 534400 633218 534458 633454
rect 534694 633218 534778 633454
rect 535014 633218 535072 633454
rect 534400 633134 535072 633218
rect 534400 632898 534458 633134
rect 534694 632898 534778 633134
rect 535014 632898 535072 633134
rect 534400 632866 535072 632898
rect 561600 633454 562272 633486
rect 561600 633218 561658 633454
rect 561894 633218 561978 633454
rect 562214 633218 562272 633454
rect 561600 633134 562272 633218
rect 561600 632898 561658 633134
rect 561894 632898 561978 633134
rect 562214 632898 562272 633134
rect 561600 632866 562272 632898
rect 571500 633454 572120 633486
rect 571500 633218 571532 633454
rect 571768 633218 571852 633454
rect 572088 633218 572120 633454
rect 571500 633134 572120 633218
rect 571500 632898 571532 633134
rect 571768 632898 571852 633134
rect 572088 632898 572120 633134
rect 571500 632866 572120 632898
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect 9084 615454 9704 615486
rect 9084 615218 9116 615454
rect 9352 615218 9436 615454
rect 9672 615218 9704 615454
rect 9084 615134 9704 615218
rect 9084 614898 9116 615134
rect 9352 614898 9436 615134
rect 9672 614898 9704 615134
rect 9084 614866 9704 614898
rect 31200 615454 31872 615486
rect 31200 615218 31258 615454
rect 31494 615218 31578 615454
rect 31814 615218 31872 615454
rect 31200 615134 31872 615218
rect 31200 614898 31258 615134
rect 31494 614898 31578 615134
rect 31814 614898 31872 615134
rect 31200 614866 31872 614898
rect 58400 615454 59072 615486
rect 58400 615218 58458 615454
rect 58694 615218 58778 615454
rect 59014 615218 59072 615454
rect 58400 615134 59072 615218
rect 58400 614898 58458 615134
rect 58694 614898 58778 615134
rect 59014 614898 59072 615134
rect 58400 614866 59072 614898
rect 85600 615454 86272 615486
rect 85600 615218 85658 615454
rect 85894 615218 85978 615454
rect 86214 615218 86272 615454
rect 85600 615134 86272 615218
rect 85600 614898 85658 615134
rect 85894 614898 85978 615134
rect 86214 614898 86272 615134
rect 85600 614866 86272 614898
rect 112800 615454 113472 615486
rect 112800 615218 112858 615454
rect 113094 615218 113178 615454
rect 113414 615218 113472 615454
rect 112800 615134 113472 615218
rect 112800 614898 112858 615134
rect 113094 614898 113178 615134
rect 113414 614898 113472 615134
rect 112800 614866 113472 614898
rect 140000 615454 140672 615486
rect 140000 615218 140058 615454
rect 140294 615218 140378 615454
rect 140614 615218 140672 615454
rect 140000 615134 140672 615218
rect 140000 614898 140058 615134
rect 140294 614898 140378 615134
rect 140614 614898 140672 615134
rect 140000 614866 140672 614898
rect 167200 615454 167872 615486
rect 167200 615218 167258 615454
rect 167494 615218 167578 615454
rect 167814 615218 167872 615454
rect 167200 615134 167872 615218
rect 167200 614898 167258 615134
rect 167494 614898 167578 615134
rect 167814 614898 167872 615134
rect 167200 614866 167872 614898
rect 194400 615454 195072 615486
rect 194400 615218 194458 615454
rect 194694 615218 194778 615454
rect 195014 615218 195072 615454
rect 194400 615134 195072 615218
rect 194400 614898 194458 615134
rect 194694 614898 194778 615134
rect 195014 614898 195072 615134
rect 194400 614866 195072 614898
rect 221600 615454 222272 615486
rect 221600 615218 221658 615454
rect 221894 615218 221978 615454
rect 222214 615218 222272 615454
rect 221600 615134 222272 615218
rect 221600 614898 221658 615134
rect 221894 614898 221978 615134
rect 222214 614898 222272 615134
rect 221600 614866 222272 614898
rect 248800 615454 249472 615486
rect 248800 615218 248858 615454
rect 249094 615218 249178 615454
rect 249414 615218 249472 615454
rect 248800 615134 249472 615218
rect 248800 614898 248858 615134
rect 249094 614898 249178 615134
rect 249414 614898 249472 615134
rect 248800 614866 249472 614898
rect 276000 615454 276672 615486
rect 276000 615218 276058 615454
rect 276294 615218 276378 615454
rect 276614 615218 276672 615454
rect 276000 615134 276672 615218
rect 276000 614898 276058 615134
rect 276294 614898 276378 615134
rect 276614 614898 276672 615134
rect 276000 614866 276672 614898
rect 303200 615454 303872 615486
rect 303200 615218 303258 615454
rect 303494 615218 303578 615454
rect 303814 615218 303872 615454
rect 303200 615134 303872 615218
rect 303200 614898 303258 615134
rect 303494 614898 303578 615134
rect 303814 614898 303872 615134
rect 303200 614866 303872 614898
rect 330400 615454 331072 615486
rect 330400 615218 330458 615454
rect 330694 615218 330778 615454
rect 331014 615218 331072 615454
rect 330400 615134 331072 615218
rect 330400 614898 330458 615134
rect 330694 614898 330778 615134
rect 331014 614898 331072 615134
rect 330400 614866 331072 614898
rect 357600 615454 358272 615486
rect 357600 615218 357658 615454
rect 357894 615218 357978 615454
rect 358214 615218 358272 615454
rect 357600 615134 358272 615218
rect 357600 614898 357658 615134
rect 357894 614898 357978 615134
rect 358214 614898 358272 615134
rect 357600 614866 358272 614898
rect 384800 615454 385472 615486
rect 384800 615218 384858 615454
rect 385094 615218 385178 615454
rect 385414 615218 385472 615454
rect 384800 615134 385472 615218
rect 384800 614898 384858 615134
rect 385094 614898 385178 615134
rect 385414 614898 385472 615134
rect 384800 614866 385472 614898
rect 412000 615454 412672 615486
rect 412000 615218 412058 615454
rect 412294 615218 412378 615454
rect 412614 615218 412672 615454
rect 412000 615134 412672 615218
rect 412000 614898 412058 615134
rect 412294 614898 412378 615134
rect 412614 614898 412672 615134
rect 412000 614866 412672 614898
rect 439200 615454 439872 615486
rect 439200 615218 439258 615454
rect 439494 615218 439578 615454
rect 439814 615218 439872 615454
rect 439200 615134 439872 615218
rect 439200 614898 439258 615134
rect 439494 614898 439578 615134
rect 439814 614898 439872 615134
rect 439200 614866 439872 614898
rect 466400 615454 467072 615486
rect 466400 615218 466458 615454
rect 466694 615218 466778 615454
rect 467014 615218 467072 615454
rect 466400 615134 467072 615218
rect 466400 614898 466458 615134
rect 466694 614898 466778 615134
rect 467014 614898 467072 615134
rect 466400 614866 467072 614898
rect 493600 615454 494272 615486
rect 493600 615218 493658 615454
rect 493894 615218 493978 615454
rect 494214 615218 494272 615454
rect 493600 615134 494272 615218
rect 493600 614898 493658 615134
rect 493894 614898 493978 615134
rect 494214 614898 494272 615134
rect 493600 614866 494272 614898
rect 520800 615454 521472 615486
rect 520800 615218 520858 615454
rect 521094 615218 521178 615454
rect 521414 615218 521472 615454
rect 520800 615134 521472 615218
rect 520800 614898 520858 615134
rect 521094 614898 521178 615134
rect 521414 614898 521472 615134
rect 520800 614866 521472 614898
rect 548000 615454 548672 615486
rect 548000 615218 548058 615454
rect 548294 615218 548378 615454
rect 548614 615218 548672 615454
rect 548000 615134 548672 615218
rect 548000 614898 548058 615134
rect 548294 614898 548378 615134
rect 548614 614898 548672 615134
rect 548000 614866 548672 614898
rect 570260 615454 570880 615486
rect 570260 615218 570292 615454
rect 570528 615218 570612 615454
rect 570848 615218 570880 615454
rect 570260 615134 570880 615218
rect 570260 614898 570292 615134
rect 570528 614898 570612 615134
rect 570848 614898 570880 615134
rect 570260 614866 570880 614898
rect 7844 597454 8464 597486
rect 7844 597218 7876 597454
rect 8112 597218 8196 597454
rect 8432 597218 8464 597454
rect 7844 597134 8464 597218
rect 7844 596898 7876 597134
rect 8112 596898 8196 597134
rect 8432 596898 8464 597134
rect 7844 596866 8464 596898
rect 17600 597454 18272 597486
rect 17600 597218 17658 597454
rect 17894 597218 17978 597454
rect 18214 597218 18272 597454
rect 17600 597134 18272 597218
rect 17600 596898 17658 597134
rect 17894 596898 17978 597134
rect 18214 596898 18272 597134
rect 17600 596866 18272 596898
rect 34835 597454 35195 597486
rect 34835 597218 34897 597454
rect 35133 597218 35195 597454
rect 34835 597134 35195 597218
rect 34835 596898 34897 597134
rect 35133 596898 35195 597134
rect 34835 596866 35195 596898
rect 133311 597454 133671 597486
rect 133311 597218 133373 597454
rect 133609 597218 133671 597454
rect 133311 597134 133671 597218
rect 133311 596898 133373 597134
rect 133609 596898 133671 597134
rect 133311 596866 133671 596898
rect 138807 597454 139167 597486
rect 138807 597218 138869 597454
rect 139105 597218 139167 597454
rect 138807 597134 139167 597218
rect 138807 596898 138869 597134
rect 139105 596898 139167 597134
rect 138807 596866 139167 596898
rect 237283 597454 237643 597486
rect 237283 597218 237345 597454
rect 237581 597218 237643 597454
rect 237283 597134 237643 597218
rect 237283 596898 237345 597134
rect 237581 596898 237643 597134
rect 237283 596866 237643 596898
rect 262400 597454 263072 597486
rect 262400 597218 262458 597454
rect 262694 597218 262778 597454
rect 263014 597218 263072 597454
rect 262400 597134 263072 597218
rect 262400 596898 262458 597134
rect 262694 596898 262778 597134
rect 263014 596898 263072 597134
rect 262400 596866 263072 596898
rect 289600 597454 290272 597486
rect 289600 597218 289658 597454
rect 289894 597218 289978 597454
rect 290214 597218 290272 597454
rect 289600 597134 290272 597218
rect 289600 596898 289658 597134
rect 289894 596898 289978 597134
rect 290214 596898 290272 597134
rect 289600 596866 290272 596898
rect 316800 597454 317472 597486
rect 316800 597218 316858 597454
rect 317094 597218 317178 597454
rect 317414 597218 317472 597454
rect 316800 597134 317472 597218
rect 316800 596898 316858 597134
rect 317094 596898 317178 597134
rect 317414 596898 317472 597134
rect 316800 596866 317472 596898
rect 341763 597454 342123 597486
rect 341763 597218 341825 597454
rect 342061 597218 342123 597454
rect 341763 597134 342123 597218
rect 341763 596898 341825 597134
rect 342061 596898 342123 597134
rect 341763 596866 342123 596898
rect 440239 597454 440599 597486
rect 440239 597218 440301 597454
rect 440537 597218 440599 597454
rect 440239 597134 440599 597218
rect 440239 596898 440301 597134
rect 440537 596898 440599 597134
rect 440239 596866 440599 596898
rect 445735 597454 446095 597486
rect 445735 597218 445797 597454
rect 446033 597218 446095 597454
rect 445735 597134 446095 597218
rect 445735 596898 445797 597134
rect 446033 596898 446095 597134
rect 445735 596866 446095 596898
rect 544211 597454 544571 597486
rect 544211 597218 544273 597454
rect 544509 597218 544571 597454
rect 544211 597134 544571 597218
rect 544211 596898 544273 597134
rect 544509 596898 544571 597134
rect 544211 596866 544571 596898
rect 561600 597454 562272 597486
rect 561600 597218 561658 597454
rect 561894 597218 561978 597454
rect 562214 597218 562272 597454
rect 561600 597134 562272 597218
rect 561600 596898 561658 597134
rect 561894 596898 561978 597134
rect 562214 596898 562272 597134
rect 561600 596866 562272 596898
rect 571500 597454 572120 597486
rect 571500 597218 571532 597454
rect 571768 597218 571852 597454
rect 572088 597218 572120 597454
rect 571500 597134 572120 597218
rect 571500 596898 571532 597134
rect 571768 596898 571852 597134
rect 572088 596898 572120 597134
rect 571500 596866 572120 596898
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect 9084 579454 9704 579486
rect 9084 579218 9116 579454
rect 9352 579218 9436 579454
rect 9672 579218 9704 579454
rect 9084 579134 9704 579218
rect 9084 578898 9116 579134
rect 9352 578898 9436 579134
rect 9672 578898 9704 579134
rect 9084 578866 9704 578898
rect 31200 579454 31872 579486
rect 31200 579218 31258 579454
rect 31494 579218 31578 579454
rect 31814 579218 31872 579454
rect 31200 579134 31872 579218
rect 31200 578898 31258 579134
rect 31494 578898 31578 579134
rect 31814 578898 31872 579134
rect 31200 578866 31872 578898
rect 35555 579454 35915 579486
rect 35555 579218 35617 579454
rect 35853 579218 35915 579454
rect 35555 579134 35915 579218
rect 35555 578898 35617 579134
rect 35853 578898 35915 579134
rect 35555 578866 35915 578898
rect 132591 579454 132951 579486
rect 132591 579218 132653 579454
rect 132889 579218 132951 579454
rect 132591 579134 132951 579218
rect 132591 578898 132653 579134
rect 132889 578898 132951 579134
rect 132591 578866 132951 578898
rect 139527 579454 139887 579486
rect 139527 579218 139589 579454
rect 139825 579218 139887 579454
rect 139527 579134 139887 579218
rect 139527 578898 139589 579134
rect 139825 578898 139887 579134
rect 139527 578866 139887 578898
rect 236563 579454 236923 579486
rect 236563 579218 236625 579454
rect 236861 579218 236923 579454
rect 236563 579134 236923 579218
rect 236563 578898 236625 579134
rect 236861 578898 236923 579134
rect 236563 578866 236923 578898
rect 248800 579454 249472 579486
rect 248800 579218 248858 579454
rect 249094 579218 249178 579454
rect 249414 579218 249472 579454
rect 248800 579134 249472 579218
rect 248800 578898 248858 579134
rect 249094 578898 249178 579134
rect 249414 578898 249472 579134
rect 248800 578866 249472 578898
rect 276000 579454 276672 579486
rect 276000 579218 276058 579454
rect 276294 579218 276378 579454
rect 276614 579218 276672 579454
rect 276000 579134 276672 579218
rect 276000 578898 276058 579134
rect 276294 578898 276378 579134
rect 276614 578898 276672 579134
rect 276000 578866 276672 578898
rect 303200 579454 303872 579486
rect 303200 579218 303258 579454
rect 303494 579218 303578 579454
rect 303814 579218 303872 579454
rect 303200 579134 303872 579218
rect 303200 578898 303258 579134
rect 303494 578898 303578 579134
rect 303814 578898 303872 579134
rect 303200 578866 303872 578898
rect 330400 579454 331072 579486
rect 330400 579218 330458 579454
rect 330694 579218 330778 579454
rect 331014 579218 331072 579454
rect 330400 579134 331072 579218
rect 330400 578898 330458 579134
rect 330694 578898 330778 579134
rect 331014 578898 331072 579134
rect 330400 578866 331072 578898
rect 342483 579454 342843 579486
rect 342483 579218 342545 579454
rect 342781 579218 342843 579454
rect 342483 579134 342843 579218
rect 342483 578898 342545 579134
rect 342781 578898 342843 579134
rect 342483 578866 342843 578898
rect 439519 579454 439879 579486
rect 439519 579218 439581 579454
rect 439817 579218 439879 579454
rect 439519 579134 439879 579218
rect 439519 578898 439581 579134
rect 439817 578898 439879 579134
rect 439519 578866 439879 578898
rect 446455 579454 446815 579486
rect 446455 579218 446517 579454
rect 446753 579218 446815 579454
rect 446455 579134 446815 579218
rect 446455 578898 446517 579134
rect 446753 578898 446815 579134
rect 446455 578866 446815 578898
rect 543491 579454 543851 579486
rect 543491 579218 543553 579454
rect 543789 579218 543851 579454
rect 543491 579134 543851 579218
rect 543491 578898 543553 579134
rect 543789 578898 543851 579134
rect 543491 578866 543851 578898
rect 548000 579454 548672 579486
rect 548000 579218 548058 579454
rect 548294 579218 548378 579454
rect 548614 579218 548672 579454
rect 548000 579134 548672 579218
rect 548000 578898 548058 579134
rect 548294 578898 548378 579134
rect 548614 578898 548672 579134
rect 548000 578866 548672 578898
rect 570260 579454 570880 579486
rect 570260 579218 570292 579454
rect 570528 579218 570612 579454
rect 570848 579218 570880 579454
rect 570260 579134 570880 579218
rect 570260 578898 570292 579134
rect 570528 578898 570612 579134
rect 570848 578898 570880 579134
rect 570260 578866 570880 578898
rect 7844 561454 8464 561486
rect 7844 561218 7876 561454
rect 8112 561218 8196 561454
rect 8432 561218 8464 561454
rect 7844 561134 8464 561218
rect 7844 560898 7876 561134
rect 8112 560898 8196 561134
rect 8432 560898 8464 561134
rect 7844 560866 8464 560898
rect 17600 561454 18272 561486
rect 17600 561218 17658 561454
rect 17894 561218 17978 561454
rect 18214 561218 18272 561454
rect 17600 561134 18272 561218
rect 17600 560898 17658 561134
rect 17894 560898 17978 561134
rect 18214 560898 18272 561134
rect 17600 560866 18272 560898
rect 34835 561454 35195 561486
rect 34835 561218 34897 561454
rect 35133 561218 35195 561454
rect 34835 561134 35195 561218
rect 34835 560898 34897 561134
rect 35133 560898 35195 561134
rect 34835 560866 35195 560898
rect 133311 561454 133671 561486
rect 133311 561218 133373 561454
rect 133609 561218 133671 561454
rect 133311 561134 133671 561218
rect 133311 560898 133373 561134
rect 133609 560898 133671 561134
rect 133311 560866 133671 560898
rect 138807 561454 139167 561486
rect 138807 561218 138869 561454
rect 139105 561218 139167 561454
rect 138807 561134 139167 561218
rect 138807 560898 138869 561134
rect 139105 560898 139167 561134
rect 138807 560866 139167 560898
rect 237283 561454 237643 561486
rect 237283 561218 237345 561454
rect 237581 561218 237643 561454
rect 237283 561134 237643 561218
rect 237283 560898 237345 561134
rect 237581 560898 237643 561134
rect 237283 560866 237643 560898
rect 262400 561454 263072 561486
rect 262400 561218 262458 561454
rect 262694 561218 262778 561454
rect 263014 561218 263072 561454
rect 262400 561134 263072 561218
rect 262400 560898 262458 561134
rect 262694 560898 262778 561134
rect 263014 560898 263072 561134
rect 262400 560866 263072 560898
rect 289600 561454 290272 561486
rect 289600 561218 289658 561454
rect 289894 561218 289978 561454
rect 290214 561218 290272 561454
rect 289600 561134 290272 561218
rect 289600 560898 289658 561134
rect 289894 560898 289978 561134
rect 290214 560898 290272 561134
rect 289600 560866 290272 560898
rect 316800 561454 317472 561486
rect 316800 561218 316858 561454
rect 317094 561218 317178 561454
rect 317414 561218 317472 561454
rect 316800 561134 317472 561218
rect 316800 560898 316858 561134
rect 317094 560898 317178 561134
rect 317414 560898 317472 561134
rect 316800 560866 317472 560898
rect 341763 561454 342123 561486
rect 341763 561218 341825 561454
rect 342061 561218 342123 561454
rect 341763 561134 342123 561218
rect 341763 560898 341825 561134
rect 342061 560898 342123 561134
rect 341763 560866 342123 560898
rect 440239 561454 440599 561486
rect 440239 561218 440301 561454
rect 440537 561218 440599 561454
rect 440239 561134 440599 561218
rect 440239 560898 440301 561134
rect 440537 560898 440599 561134
rect 440239 560866 440599 560898
rect 445735 561454 446095 561486
rect 445735 561218 445797 561454
rect 446033 561218 446095 561454
rect 445735 561134 446095 561218
rect 445735 560898 445797 561134
rect 446033 560898 446095 561134
rect 445735 560866 446095 560898
rect 544211 561454 544571 561486
rect 544211 561218 544273 561454
rect 544509 561218 544571 561454
rect 544211 561134 544571 561218
rect 544211 560898 544273 561134
rect 544509 560898 544571 561134
rect 544211 560866 544571 560898
rect 561600 561454 562272 561486
rect 561600 561218 561658 561454
rect 561894 561218 561978 561454
rect 562214 561218 562272 561454
rect 561600 561134 562272 561218
rect 561600 560898 561658 561134
rect 561894 560898 561978 561134
rect 562214 560898 562272 561134
rect 561600 560866 562272 560898
rect 571500 561454 572120 561486
rect 571500 561218 571532 561454
rect 571768 561218 571852 561454
rect 572088 561218 572120 561454
rect 571500 561134 572120 561218
rect 571500 560898 571532 561134
rect 571768 560898 571852 561134
rect 572088 560898 572120 561134
rect 571500 560866 572120 560898
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect 9084 543454 9704 543486
rect 9084 543218 9116 543454
rect 9352 543218 9436 543454
rect 9672 543218 9704 543454
rect 9084 543134 9704 543218
rect 9084 542898 9116 543134
rect 9352 542898 9436 543134
rect 9672 542898 9704 543134
rect 9084 542866 9704 542898
rect 31200 543454 31872 543486
rect 31200 543218 31258 543454
rect 31494 543218 31578 543454
rect 31814 543218 31872 543454
rect 31200 543134 31872 543218
rect 31200 542898 31258 543134
rect 31494 542898 31578 543134
rect 31814 542898 31872 543134
rect 31200 542866 31872 542898
rect 35555 543454 35915 543486
rect 35555 543218 35617 543454
rect 35853 543218 35915 543454
rect 35555 543134 35915 543218
rect 35555 542898 35617 543134
rect 35853 542898 35915 543134
rect 35555 542866 35915 542898
rect 132591 543454 132951 543486
rect 132591 543218 132653 543454
rect 132889 543218 132951 543454
rect 132591 543134 132951 543218
rect 132591 542898 132653 543134
rect 132889 542898 132951 543134
rect 132591 542866 132951 542898
rect 139527 543454 139887 543486
rect 139527 543218 139589 543454
rect 139825 543218 139887 543454
rect 139527 543134 139887 543218
rect 139527 542898 139589 543134
rect 139825 542898 139887 543134
rect 139527 542866 139887 542898
rect 236563 543454 236923 543486
rect 236563 543218 236625 543454
rect 236861 543218 236923 543454
rect 236563 543134 236923 543218
rect 236563 542898 236625 543134
rect 236861 542898 236923 543134
rect 236563 542866 236923 542898
rect 248800 543454 249472 543486
rect 248800 543218 248858 543454
rect 249094 543218 249178 543454
rect 249414 543218 249472 543454
rect 248800 543134 249472 543218
rect 248800 542898 248858 543134
rect 249094 542898 249178 543134
rect 249414 542898 249472 543134
rect 248800 542866 249472 542898
rect 276000 543454 276672 543486
rect 276000 543218 276058 543454
rect 276294 543218 276378 543454
rect 276614 543218 276672 543454
rect 276000 543134 276672 543218
rect 276000 542898 276058 543134
rect 276294 542898 276378 543134
rect 276614 542898 276672 543134
rect 276000 542866 276672 542898
rect 303200 543454 303872 543486
rect 303200 543218 303258 543454
rect 303494 543218 303578 543454
rect 303814 543218 303872 543454
rect 303200 543134 303872 543218
rect 303200 542898 303258 543134
rect 303494 542898 303578 543134
rect 303814 542898 303872 543134
rect 303200 542866 303872 542898
rect 330400 543454 331072 543486
rect 330400 543218 330458 543454
rect 330694 543218 330778 543454
rect 331014 543218 331072 543454
rect 330400 543134 331072 543218
rect 330400 542898 330458 543134
rect 330694 542898 330778 543134
rect 331014 542898 331072 543134
rect 330400 542866 331072 542898
rect 342483 543454 342843 543486
rect 342483 543218 342545 543454
rect 342781 543218 342843 543454
rect 342483 543134 342843 543218
rect 342483 542898 342545 543134
rect 342781 542898 342843 543134
rect 342483 542866 342843 542898
rect 439519 543454 439879 543486
rect 439519 543218 439581 543454
rect 439817 543218 439879 543454
rect 439519 543134 439879 543218
rect 439519 542898 439581 543134
rect 439817 542898 439879 543134
rect 439519 542866 439879 542898
rect 446455 543454 446815 543486
rect 446455 543218 446517 543454
rect 446753 543218 446815 543454
rect 446455 543134 446815 543218
rect 446455 542898 446517 543134
rect 446753 542898 446815 543134
rect 446455 542866 446815 542898
rect 543491 543454 543851 543486
rect 543491 543218 543553 543454
rect 543789 543218 543851 543454
rect 543491 543134 543851 543218
rect 543491 542898 543553 543134
rect 543789 542898 543851 543134
rect 543491 542866 543851 542898
rect 548000 543454 548672 543486
rect 548000 543218 548058 543454
rect 548294 543218 548378 543454
rect 548614 543218 548672 543454
rect 548000 543134 548672 543218
rect 548000 542898 548058 543134
rect 548294 542898 548378 543134
rect 548614 542898 548672 543134
rect 548000 542866 548672 542898
rect 570260 543454 570880 543486
rect 570260 543218 570292 543454
rect 570528 543218 570612 543454
rect 570848 543218 570880 543454
rect 570260 543134 570880 543218
rect 570260 542898 570292 543134
rect 570528 542898 570612 543134
rect 570848 542898 570880 543134
rect 570260 542866 570880 542898
rect 7844 525454 8464 525486
rect 7844 525218 7876 525454
rect 8112 525218 8196 525454
rect 8432 525218 8464 525454
rect 7844 525134 8464 525218
rect 7844 524898 7876 525134
rect 8112 524898 8196 525134
rect 8432 524898 8464 525134
rect 7844 524866 8464 524898
rect 17600 525454 18272 525486
rect 17600 525218 17658 525454
rect 17894 525218 17978 525454
rect 18214 525218 18272 525454
rect 17600 525134 18272 525218
rect 17600 524898 17658 525134
rect 17894 524898 17978 525134
rect 18214 524898 18272 525134
rect 17600 524866 18272 524898
rect 44800 525454 45472 525486
rect 44800 525218 44858 525454
rect 45094 525218 45178 525454
rect 45414 525218 45472 525454
rect 44800 525134 45472 525218
rect 44800 524898 44858 525134
rect 45094 524898 45178 525134
rect 45414 524898 45472 525134
rect 44800 524866 45472 524898
rect 72000 525454 72672 525486
rect 72000 525218 72058 525454
rect 72294 525218 72378 525454
rect 72614 525218 72672 525454
rect 72000 525134 72672 525218
rect 72000 524898 72058 525134
rect 72294 524898 72378 525134
rect 72614 524898 72672 525134
rect 72000 524866 72672 524898
rect 99200 525454 99872 525486
rect 99200 525218 99258 525454
rect 99494 525218 99578 525454
rect 99814 525218 99872 525454
rect 99200 525134 99872 525218
rect 99200 524898 99258 525134
rect 99494 524898 99578 525134
rect 99814 524898 99872 525134
rect 99200 524866 99872 524898
rect 126400 525454 127072 525486
rect 126400 525218 126458 525454
rect 126694 525218 126778 525454
rect 127014 525218 127072 525454
rect 126400 525134 127072 525218
rect 126400 524898 126458 525134
rect 126694 524898 126778 525134
rect 127014 524898 127072 525134
rect 126400 524866 127072 524898
rect 153600 525454 154272 525486
rect 153600 525218 153658 525454
rect 153894 525218 153978 525454
rect 154214 525218 154272 525454
rect 153600 525134 154272 525218
rect 153600 524898 153658 525134
rect 153894 524898 153978 525134
rect 154214 524898 154272 525134
rect 153600 524866 154272 524898
rect 180800 525454 181472 525486
rect 180800 525218 180858 525454
rect 181094 525218 181178 525454
rect 181414 525218 181472 525454
rect 180800 525134 181472 525218
rect 180800 524898 180858 525134
rect 181094 524898 181178 525134
rect 181414 524898 181472 525134
rect 180800 524866 181472 524898
rect 208000 525454 208672 525486
rect 208000 525218 208058 525454
rect 208294 525218 208378 525454
rect 208614 525218 208672 525454
rect 208000 525134 208672 525218
rect 208000 524898 208058 525134
rect 208294 524898 208378 525134
rect 208614 524898 208672 525134
rect 208000 524866 208672 524898
rect 235200 525454 235872 525486
rect 235200 525218 235258 525454
rect 235494 525218 235578 525454
rect 235814 525218 235872 525454
rect 235200 525134 235872 525218
rect 235200 524898 235258 525134
rect 235494 524898 235578 525134
rect 235814 524898 235872 525134
rect 235200 524866 235872 524898
rect 262400 525454 263072 525486
rect 262400 525218 262458 525454
rect 262694 525218 262778 525454
rect 263014 525218 263072 525454
rect 262400 525134 263072 525218
rect 262400 524898 262458 525134
rect 262694 524898 262778 525134
rect 263014 524898 263072 525134
rect 262400 524866 263072 524898
rect 289600 525454 290272 525486
rect 289600 525218 289658 525454
rect 289894 525218 289978 525454
rect 290214 525218 290272 525454
rect 289600 525134 290272 525218
rect 289600 524898 289658 525134
rect 289894 524898 289978 525134
rect 290214 524898 290272 525134
rect 289600 524866 290272 524898
rect 316800 525454 317472 525486
rect 316800 525218 316858 525454
rect 317094 525218 317178 525454
rect 317414 525218 317472 525454
rect 316800 525134 317472 525218
rect 316800 524898 316858 525134
rect 317094 524898 317178 525134
rect 317414 524898 317472 525134
rect 316800 524866 317472 524898
rect 344000 525454 344672 525486
rect 344000 525218 344058 525454
rect 344294 525218 344378 525454
rect 344614 525218 344672 525454
rect 344000 525134 344672 525218
rect 344000 524898 344058 525134
rect 344294 524898 344378 525134
rect 344614 524898 344672 525134
rect 344000 524866 344672 524898
rect 371200 525454 371872 525486
rect 371200 525218 371258 525454
rect 371494 525218 371578 525454
rect 371814 525218 371872 525454
rect 371200 525134 371872 525218
rect 371200 524898 371258 525134
rect 371494 524898 371578 525134
rect 371814 524898 371872 525134
rect 371200 524866 371872 524898
rect 398400 525454 399072 525486
rect 398400 525218 398458 525454
rect 398694 525218 398778 525454
rect 399014 525218 399072 525454
rect 398400 525134 399072 525218
rect 398400 524898 398458 525134
rect 398694 524898 398778 525134
rect 399014 524898 399072 525134
rect 398400 524866 399072 524898
rect 425600 525454 426272 525486
rect 425600 525218 425658 525454
rect 425894 525218 425978 525454
rect 426214 525218 426272 525454
rect 425600 525134 426272 525218
rect 425600 524898 425658 525134
rect 425894 524898 425978 525134
rect 426214 524898 426272 525134
rect 425600 524866 426272 524898
rect 452800 525454 453472 525486
rect 452800 525218 452858 525454
rect 453094 525218 453178 525454
rect 453414 525218 453472 525454
rect 452800 525134 453472 525218
rect 452800 524898 452858 525134
rect 453094 524898 453178 525134
rect 453414 524898 453472 525134
rect 452800 524866 453472 524898
rect 480000 525454 480672 525486
rect 480000 525218 480058 525454
rect 480294 525218 480378 525454
rect 480614 525218 480672 525454
rect 480000 525134 480672 525218
rect 480000 524898 480058 525134
rect 480294 524898 480378 525134
rect 480614 524898 480672 525134
rect 480000 524866 480672 524898
rect 507200 525454 507872 525486
rect 507200 525218 507258 525454
rect 507494 525218 507578 525454
rect 507814 525218 507872 525454
rect 507200 525134 507872 525218
rect 507200 524898 507258 525134
rect 507494 524898 507578 525134
rect 507814 524898 507872 525134
rect 507200 524866 507872 524898
rect 534400 525454 535072 525486
rect 534400 525218 534458 525454
rect 534694 525218 534778 525454
rect 535014 525218 535072 525454
rect 534400 525134 535072 525218
rect 534400 524898 534458 525134
rect 534694 524898 534778 525134
rect 535014 524898 535072 525134
rect 534400 524866 535072 524898
rect 561600 525454 562272 525486
rect 561600 525218 561658 525454
rect 561894 525218 561978 525454
rect 562214 525218 562272 525454
rect 561600 525134 562272 525218
rect 561600 524898 561658 525134
rect 561894 524898 561978 525134
rect 562214 524898 562272 525134
rect 561600 524866 562272 524898
rect 571500 525454 572120 525486
rect 571500 525218 571532 525454
rect 571768 525218 571852 525454
rect 572088 525218 572120 525454
rect 571500 525134 572120 525218
rect 571500 524898 571532 525134
rect 571768 524898 571852 525134
rect 572088 524898 572120 525134
rect 571500 524866 572120 524898
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect 9084 507454 9704 507486
rect 9084 507218 9116 507454
rect 9352 507218 9436 507454
rect 9672 507218 9704 507454
rect 9084 507134 9704 507218
rect 9084 506898 9116 507134
rect 9352 506898 9436 507134
rect 9672 506898 9704 507134
rect 9084 506866 9704 506898
rect 31200 507454 31872 507486
rect 31200 507218 31258 507454
rect 31494 507218 31578 507454
rect 31814 507218 31872 507454
rect 31200 507134 31872 507218
rect 31200 506898 31258 507134
rect 31494 506898 31578 507134
rect 31814 506898 31872 507134
rect 31200 506866 31872 506898
rect 35555 507454 35915 507486
rect 35555 507218 35617 507454
rect 35853 507218 35915 507454
rect 35555 507134 35915 507218
rect 35555 506898 35617 507134
rect 35853 506898 35915 507134
rect 35555 506866 35915 506898
rect 132591 507454 132951 507486
rect 132591 507218 132653 507454
rect 132889 507218 132951 507454
rect 132591 507134 132951 507218
rect 132591 506898 132653 507134
rect 132889 506898 132951 507134
rect 132591 506866 132951 506898
rect 139527 507454 139887 507486
rect 139527 507218 139589 507454
rect 139825 507218 139887 507454
rect 139527 507134 139887 507218
rect 139527 506898 139589 507134
rect 139825 506898 139887 507134
rect 139527 506866 139887 506898
rect 236563 507454 236923 507486
rect 236563 507218 236625 507454
rect 236861 507218 236923 507454
rect 236563 507134 236923 507218
rect 236563 506898 236625 507134
rect 236861 506898 236923 507134
rect 236563 506866 236923 506898
rect 248800 507454 249472 507486
rect 248800 507218 248858 507454
rect 249094 507218 249178 507454
rect 249414 507218 249472 507454
rect 248800 507134 249472 507218
rect 248800 506898 248858 507134
rect 249094 506898 249178 507134
rect 249414 506898 249472 507134
rect 248800 506866 249472 506898
rect 276000 507454 276672 507486
rect 276000 507218 276058 507454
rect 276294 507218 276378 507454
rect 276614 507218 276672 507454
rect 276000 507134 276672 507218
rect 276000 506898 276058 507134
rect 276294 506898 276378 507134
rect 276614 506898 276672 507134
rect 276000 506866 276672 506898
rect 303200 507454 303872 507486
rect 303200 507218 303258 507454
rect 303494 507218 303578 507454
rect 303814 507218 303872 507454
rect 303200 507134 303872 507218
rect 303200 506898 303258 507134
rect 303494 506898 303578 507134
rect 303814 506898 303872 507134
rect 303200 506866 303872 506898
rect 330400 507454 331072 507486
rect 330400 507218 330458 507454
rect 330694 507218 330778 507454
rect 331014 507218 331072 507454
rect 330400 507134 331072 507218
rect 330400 506898 330458 507134
rect 330694 506898 330778 507134
rect 331014 506898 331072 507134
rect 330400 506866 331072 506898
rect 342483 507454 342843 507486
rect 342483 507218 342545 507454
rect 342781 507218 342843 507454
rect 342483 507134 342843 507218
rect 342483 506898 342545 507134
rect 342781 506898 342843 507134
rect 342483 506866 342843 506898
rect 439519 507454 439879 507486
rect 439519 507218 439581 507454
rect 439817 507218 439879 507454
rect 439519 507134 439879 507218
rect 439519 506898 439581 507134
rect 439817 506898 439879 507134
rect 439519 506866 439879 506898
rect 446455 507454 446815 507486
rect 446455 507218 446517 507454
rect 446753 507218 446815 507454
rect 446455 507134 446815 507218
rect 446455 506898 446517 507134
rect 446753 506898 446815 507134
rect 446455 506866 446815 506898
rect 543491 507454 543851 507486
rect 543491 507218 543553 507454
rect 543789 507218 543851 507454
rect 543491 507134 543851 507218
rect 543491 506898 543553 507134
rect 543789 506898 543851 507134
rect 543491 506866 543851 506898
rect 548000 507454 548672 507486
rect 548000 507218 548058 507454
rect 548294 507218 548378 507454
rect 548614 507218 548672 507454
rect 548000 507134 548672 507218
rect 548000 506898 548058 507134
rect 548294 506898 548378 507134
rect 548614 506898 548672 507134
rect 548000 506866 548672 506898
rect 570260 507454 570880 507486
rect 570260 507218 570292 507454
rect 570528 507218 570612 507454
rect 570848 507218 570880 507454
rect 570260 507134 570880 507218
rect 570260 506898 570292 507134
rect 570528 506898 570612 507134
rect 570848 506898 570880 507134
rect 570260 506866 570880 506898
rect 7844 489454 8464 489486
rect 7844 489218 7876 489454
rect 8112 489218 8196 489454
rect 8432 489218 8464 489454
rect 7844 489134 8464 489218
rect 7844 488898 7876 489134
rect 8112 488898 8196 489134
rect 8432 488898 8464 489134
rect 7844 488866 8464 488898
rect 17600 489454 18272 489486
rect 17600 489218 17658 489454
rect 17894 489218 17978 489454
rect 18214 489218 18272 489454
rect 17600 489134 18272 489218
rect 17600 488898 17658 489134
rect 17894 488898 17978 489134
rect 18214 488898 18272 489134
rect 17600 488866 18272 488898
rect 34835 489454 35195 489486
rect 34835 489218 34897 489454
rect 35133 489218 35195 489454
rect 34835 489134 35195 489218
rect 34835 488898 34897 489134
rect 35133 488898 35195 489134
rect 34835 488866 35195 488898
rect 133311 489454 133671 489486
rect 133311 489218 133373 489454
rect 133609 489218 133671 489454
rect 133311 489134 133671 489218
rect 133311 488898 133373 489134
rect 133609 488898 133671 489134
rect 133311 488866 133671 488898
rect 138807 489454 139167 489486
rect 138807 489218 138869 489454
rect 139105 489218 139167 489454
rect 138807 489134 139167 489218
rect 138807 488898 138869 489134
rect 139105 488898 139167 489134
rect 138807 488866 139167 488898
rect 237283 489454 237643 489486
rect 237283 489218 237345 489454
rect 237581 489218 237643 489454
rect 237283 489134 237643 489218
rect 237283 488898 237345 489134
rect 237581 488898 237643 489134
rect 237283 488866 237643 488898
rect 262400 489454 263072 489486
rect 262400 489218 262458 489454
rect 262694 489218 262778 489454
rect 263014 489218 263072 489454
rect 262400 489134 263072 489218
rect 262400 488898 262458 489134
rect 262694 488898 262778 489134
rect 263014 488898 263072 489134
rect 262400 488866 263072 488898
rect 289600 489454 290272 489486
rect 289600 489218 289658 489454
rect 289894 489218 289978 489454
rect 290214 489218 290272 489454
rect 289600 489134 290272 489218
rect 289600 488898 289658 489134
rect 289894 488898 289978 489134
rect 290214 488898 290272 489134
rect 289600 488866 290272 488898
rect 316800 489454 317472 489486
rect 316800 489218 316858 489454
rect 317094 489218 317178 489454
rect 317414 489218 317472 489454
rect 316800 489134 317472 489218
rect 316800 488898 316858 489134
rect 317094 488898 317178 489134
rect 317414 488898 317472 489134
rect 316800 488866 317472 488898
rect 341763 489454 342123 489486
rect 341763 489218 341825 489454
rect 342061 489218 342123 489454
rect 341763 489134 342123 489218
rect 341763 488898 341825 489134
rect 342061 488898 342123 489134
rect 341763 488866 342123 488898
rect 440239 489454 440599 489486
rect 440239 489218 440301 489454
rect 440537 489218 440599 489454
rect 440239 489134 440599 489218
rect 440239 488898 440301 489134
rect 440537 488898 440599 489134
rect 440239 488866 440599 488898
rect 445735 489454 446095 489486
rect 445735 489218 445797 489454
rect 446033 489218 446095 489454
rect 445735 489134 446095 489218
rect 445735 488898 445797 489134
rect 446033 488898 446095 489134
rect 445735 488866 446095 488898
rect 544211 489454 544571 489486
rect 544211 489218 544273 489454
rect 544509 489218 544571 489454
rect 544211 489134 544571 489218
rect 544211 488898 544273 489134
rect 544509 488898 544571 489134
rect 544211 488866 544571 488898
rect 561600 489454 562272 489486
rect 561600 489218 561658 489454
rect 561894 489218 561978 489454
rect 562214 489218 562272 489454
rect 561600 489134 562272 489218
rect 561600 488898 561658 489134
rect 561894 488898 561978 489134
rect 562214 488898 562272 489134
rect 561600 488866 562272 488898
rect 571500 489454 572120 489486
rect 571500 489218 571532 489454
rect 571768 489218 571852 489454
rect 572088 489218 572120 489454
rect 571500 489134 572120 489218
rect 571500 488898 571532 489134
rect 571768 488898 571852 489134
rect 572088 488898 572120 489134
rect 571500 488866 572120 488898
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect 9084 471454 9704 471486
rect 9084 471218 9116 471454
rect 9352 471218 9436 471454
rect 9672 471218 9704 471454
rect 9084 471134 9704 471218
rect 9084 470898 9116 471134
rect 9352 470898 9436 471134
rect 9672 470898 9704 471134
rect 9084 470866 9704 470898
rect 31200 471454 31872 471486
rect 31200 471218 31258 471454
rect 31494 471218 31578 471454
rect 31814 471218 31872 471454
rect 31200 471134 31872 471218
rect 31200 470898 31258 471134
rect 31494 470898 31578 471134
rect 31814 470898 31872 471134
rect 31200 470866 31872 470898
rect 35555 471454 35915 471486
rect 35555 471218 35617 471454
rect 35853 471218 35915 471454
rect 35555 471134 35915 471218
rect 35555 470898 35617 471134
rect 35853 470898 35915 471134
rect 35555 470866 35915 470898
rect 132591 471454 132951 471486
rect 132591 471218 132653 471454
rect 132889 471218 132951 471454
rect 132591 471134 132951 471218
rect 132591 470898 132653 471134
rect 132889 470898 132951 471134
rect 132591 470866 132951 470898
rect 139527 471454 139887 471486
rect 139527 471218 139589 471454
rect 139825 471218 139887 471454
rect 139527 471134 139887 471218
rect 139527 470898 139589 471134
rect 139825 470898 139887 471134
rect 139527 470866 139887 470898
rect 236563 471454 236923 471486
rect 236563 471218 236625 471454
rect 236861 471218 236923 471454
rect 236563 471134 236923 471218
rect 236563 470898 236625 471134
rect 236861 470898 236923 471134
rect 236563 470866 236923 470898
rect 248800 471454 249472 471486
rect 248800 471218 248858 471454
rect 249094 471218 249178 471454
rect 249414 471218 249472 471454
rect 248800 471134 249472 471218
rect 248800 470898 248858 471134
rect 249094 470898 249178 471134
rect 249414 470898 249472 471134
rect 248800 470866 249472 470898
rect 276000 471454 276672 471486
rect 276000 471218 276058 471454
rect 276294 471218 276378 471454
rect 276614 471218 276672 471454
rect 276000 471134 276672 471218
rect 276000 470898 276058 471134
rect 276294 470898 276378 471134
rect 276614 470898 276672 471134
rect 276000 470866 276672 470898
rect 303200 471454 303872 471486
rect 303200 471218 303258 471454
rect 303494 471218 303578 471454
rect 303814 471218 303872 471454
rect 303200 471134 303872 471218
rect 303200 470898 303258 471134
rect 303494 470898 303578 471134
rect 303814 470898 303872 471134
rect 303200 470866 303872 470898
rect 330400 471454 331072 471486
rect 330400 471218 330458 471454
rect 330694 471218 330778 471454
rect 331014 471218 331072 471454
rect 330400 471134 331072 471218
rect 330400 470898 330458 471134
rect 330694 470898 330778 471134
rect 331014 470898 331072 471134
rect 330400 470866 331072 470898
rect 342483 471454 342843 471486
rect 342483 471218 342545 471454
rect 342781 471218 342843 471454
rect 342483 471134 342843 471218
rect 342483 470898 342545 471134
rect 342781 470898 342843 471134
rect 342483 470866 342843 470898
rect 439519 471454 439879 471486
rect 439519 471218 439581 471454
rect 439817 471218 439879 471454
rect 439519 471134 439879 471218
rect 439519 470898 439581 471134
rect 439817 470898 439879 471134
rect 439519 470866 439879 470898
rect 446455 471454 446815 471486
rect 446455 471218 446517 471454
rect 446753 471218 446815 471454
rect 446455 471134 446815 471218
rect 446455 470898 446517 471134
rect 446753 470898 446815 471134
rect 446455 470866 446815 470898
rect 543491 471454 543851 471486
rect 543491 471218 543553 471454
rect 543789 471218 543851 471454
rect 543491 471134 543851 471218
rect 543491 470898 543553 471134
rect 543789 470898 543851 471134
rect 543491 470866 543851 470898
rect 548000 471454 548672 471486
rect 548000 471218 548058 471454
rect 548294 471218 548378 471454
rect 548614 471218 548672 471454
rect 548000 471134 548672 471218
rect 548000 470898 548058 471134
rect 548294 470898 548378 471134
rect 548614 470898 548672 471134
rect 548000 470866 548672 470898
rect 570260 471454 570880 471486
rect 570260 471218 570292 471454
rect 570528 471218 570612 471454
rect 570848 471218 570880 471454
rect 570260 471134 570880 471218
rect 570260 470898 570292 471134
rect 570528 470898 570612 471134
rect 570848 470898 570880 471134
rect 570260 470866 570880 470898
rect 7844 453454 8464 453486
rect 7844 453218 7876 453454
rect 8112 453218 8196 453454
rect 8432 453218 8464 453454
rect 7844 453134 8464 453218
rect 7844 452898 7876 453134
rect 8112 452898 8196 453134
rect 8432 452898 8464 453134
rect 7844 452866 8464 452898
rect 17600 453454 18272 453486
rect 17600 453218 17658 453454
rect 17894 453218 17978 453454
rect 18214 453218 18272 453454
rect 17600 453134 18272 453218
rect 17600 452898 17658 453134
rect 17894 452898 17978 453134
rect 18214 452898 18272 453134
rect 17600 452866 18272 452898
rect 34835 453454 35195 453486
rect 34835 453218 34897 453454
rect 35133 453218 35195 453454
rect 34835 453134 35195 453218
rect 34835 452898 34897 453134
rect 35133 452898 35195 453134
rect 34835 452866 35195 452898
rect 133311 453454 133671 453486
rect 133311 453218 133373 453454
rect 133609 453218 133671 453454
rect 133311 453134 133671 453218
rect 133311 452898 133373 453134
rect 133609 452898 133671 453134
rect 133311 452866 133671 452898
rect 138807 453454 139167 453486
rect 138807 453218 138869 453454
rect 139105 453218 139167 453454
rect 138807 453134 139167 453218
rect 138807 452898 138869 453134
rect 139105 452898 139167 453134
rect 138807 452866 139167 452898
rect 237283 453454 237643 453486
rect 237283 453218 237345 453454
rect 237581 453218 237643 453454
rect 237283 453134 237643 453218
rect 237283 452898 237345 453134
rect 237581 452898 237643 453134
rect 237283 452866 237643 452898
rect 262400 453454 263072 453486
rect 262400 453218 262458 453454
rect 262694 453218 262778 453454
rect 263014 453218 263072 453454
rect 262400 453134 263072 453218
rect 262400 452898 262458 453134
rect 262694 452898 262778 453134
rect 263014 452898 263072 453134
rect 262400 452866 263072 452898
rect 289600 453454 290272 453486
rect 289600 453218 289658 453454
rect 289894 453218 289978 453454
rect 290214 453218 290272 453454
rect 289600 453134 290272 453218
rect 289600 452898 289658 453134
rect 289894 452898 289978 453134
rect 290214 452898 290272 453134
rect 289600 452866 290272 452898
rect 316800 453454 317472 453486
rect 316800 453218 316858 453454
rect 317094 453218 317178 453454
rect 317414 453218 317472 453454
rect 316800 453134 317472 453218
rect 316800 452898 316858 453134
rect 317094 452898 317178 453134
rect 317414 452898 317472 453134
rect 316800 452866 317472 452898
rect 341763 453454 342123 453486
rect 341763 453218 341825 453454
rect 342061 453218 342123 453454
rect 341763 453134 342123 453218
rect 341763 452898 341825 453134
rect 342061 452898 342123 453134
rect 341763 452866 342123 452898
rect 440239 453454 440599 453486
rect 440239 453218 440301 453454
rect 440537 453218 440599 453454
rect 440239 453134 440599 453218
rect 440239 452898 440301 453134
rect 440537 452898 440599 453134
rect 440239 452866 440599 452898
rect 445735 453454 446095 453486
rect 445735 453218 445797 453454
rect 446033 453218 446095 453454
rect 445735 453134 446095 453218
rect 445735 452898 445797 453134
rect 446033 452898 446095 453134
rect 445735 452866 446095 452898
rect 544211 453454 544571 453486
rect 544211 453218 544273 453454
rect 544509 453218 544571 453454
rect 544211 453134 544571 453218
rect 544211 452898 544273 453134
rect 544509 452898 544571 453134
rect 544211 452866 544571 452898
rect 561600 453454 562272 453486
rect 561600 453218 561658 453454
rect 561894 453218 561978 453454
rect 562214 453218 562272 453454
rect 561600 453134 562272 453218
rect 561600 452898 561658 453134
rect 561894 452898 561978 453134
rect 562214 452898 562272 453134
rect 561600 452866 562272 452898
rect 571500 453454 572120 453486
rect 571500 453218 571532 453454
rect 571768 453218 571852 453454
rect 572088 453218 572120 453454
rect 571500 453134 572120 453218
rect 571500 452898 571532 453134
rect 571768 452898 571852 453134
rect 572088 452898 572120 453134
rect 571500 452866 572120 452898
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect 9084 435454 9704 435486
rect 9084 435218 9116 435454
rect 9352 435218 9436 435454
rect 9672 435218 9704 435454
rect 9084 435134 9704 435218
rect 9084 434898 9116 435134
rect 9352 434898 9436 435134
rect 9672 434898 9704 435134
rect 9084 434866 9704 434898
rect 31200 435454 31872 435486
rect 31200 435218 31258 435454
rect 31494 435218 31578 435454
rect 31814 435218 31872 435454
rect 31200 435134 31872 435218
rect 31200 434898 31258 435134
rect 31494 434898 31578 435134
rect 31814 434898 31872 435134
rect 31200 434866 31872 434898
rect 58400 435454 59072 435486
rect 58400 435218 58458 435454
rect 58694 435218 58778 435454
rect 59014 435218 59072 435454
rect 58400 435134 59072 435218
rect 58400 434898 58458 435134
rect 58694 434898 58778 435134
rect 59014 434898 59072 435134
rect 58400 434866 59072 434898
rect 85600 435454 86272 435486
rect 85600 435218 85658 435454
rect 85894 435218 85978 435454
rect 86214 435218 86272 435454
rect 85600 435134 86272 435218
rect 85600 434898 85658 435134
rect 85894 434898 85978 435134
rect 86214 434898 86272 435134
rect 85600 434866 86272 434898
rect 112800 435454 113472 435486
rect 112800 435218 112858 435454
rect 113094 435218 113178 435454
rect 113414 435218 113472 435454
rect 112800 435134 113472 435218
rect 112800 434898 112858 435134
rect 113094 434898 113178 435134
rect 113414 434898 113472 435134
rect 112800 434866 113472 434898
rect 140000 435454 140672 435486
rect 140000 435218 140058 435454
rect 140294 435218 140378 435454
rect 140614 435218 140672 435454
rect 140000 435134 140672 435218
rect 140000 434898 140058 435134
rect 140294 434898 140378 435134
rect 140614 434898 140672 435134
rect 140000 434866 140672 434898
rect 167200 435454 167872 435486
rect 167200 435218 167258 435454
rect 167494 435218 167578 435454
rect 167814 435218 167872 435454
rect 167200 435134 167872 435218
rect 167200 434898 167258 435134
rect 167494 434898 167578 435134
rect 167814 434898 167872 435134
rect 167200 434866 167872 434898
rect 194400 435454 195072 435486
rect 194400 435218 194458 435454
rect 194694 435218 194778 435454
rect 195014 435218 195072 435454
rect 194400 435134 195072 435218
rect 194400 434898 194458 435134
rect 194694 434898 194778 435134
rect 195014 434898 195072 435134
rect 194400 434866 195072 434898
rect 221600 435454 222272 435486
rect 221600 435218 221658 435454
rect 221894 435218 221978 435454
rect 222214 435218 222272 435454
rect 221600 435134 222272 435218
rect 221600 434898 221658 435134
rect 221894 434898 221978 435134
rect 222214 434898 222272 435134
rect 221600 434866 222272 434898
rect 248800 435454 249472 435486
rect 248800 435218 248858 435454
rect 249094 435218 249178 435454
rect 249414 435218 249472 435454
rect 248800 435134 249472 435218
rect 248800 434898 248858 435134
rect 249094 434898 249178 435134
rect 249414 434898 249472 435134
rect 248800 434866 249472 434898
rect 276000 435454 276672 435486
rect 276000 435218 276058 435454
rect 276294 435218 276378 435454
rect 276614 435218 276672 435454
rect 276000 435134 276672 435218
rect 276000 434898 276058 435134
rect 276294 434898 276378 435134
rect 276614 434898 276672 435134
rect 276000 434866 276672 434898
rect 303200 435454 303872 435486
rect 303200 435218 303258 435454
rect 303494 435218 303578 435454
rect 303814 435218 303872 435454
rect 303200 435134 303872 435218
rect 303200 434898 303258 435134
rect 303494 434898 303578 435134
rect 303814 434898 303872 435134
rect 303200 434866 303872 434898
rect 330400 435454 331072 435486
rect 330400 435218 330458 435454
rect 330694 435218 330778 435454
rect 331014 435218 331072 435454
rect 330400 435134 331072 435218
rect 330400 434898 330458 435134
rect 330694 434898 330778 435134
rect 331014 434898 331072 435134
rect 330400 434866 331072 434898
rect 357600 435454 358272 435486
rect 357600 435218 357658 435454
rect 357894 435218 357978 435454
rect 358214 435218 358272 435454
rect 357600 435134 358272 435218
rect 357600 434898 357658 435134
rect 357894 434898 357978 435134
rect 358214 434898 358272 435134
rect 357600 434866 358272 434898
rect 384800 435454 385472 435486
rect 384800 435218 384858 435454
rect 385094 435218 385178 435454
rect 385414 435218 385472 435454
rect 384800 435134 385472 435218
rect 384800 434898 384858 435134
rect 385094 434898 385178 435134
rect 385414 434898 385472 435134
rect 384800 434866 385472 434898
rect 412000 435454 412672 435486
rect 412000 435218 412058 435454
rect 412294 435218 412378 435454
rect 412614 435218 412672 435454
rect 412000 435134 412672 435218
rect 412000 434898 412058 435134
rect 412294 434898 412378 435134
rect 412614 434898 412672 435134
rect 412000 434866 412672 434898
rect 439200 435454 439872 435486
rect 439200 435218 439258 435454
rect 439494 435218 439578 435454
rect 439814 435218 439872 435454
rect 439200 435134 439872 435218
rect 439200 434898 439258 435134
rect 439494 434898 439578 435134
rect 439814 434898 439872 435134
rect 439200 434866 439872 434898
rect 466400 435454 467072 435486
rect 466400 435218 466458 435454
rect 466694 435218 466778 435454
rect 467014 435218 467072 435454
rect 466400 435134 467072 435218
rect 466400 434898 466458 435134
rect 466694 434898 466778 435134
rect 467014 434898 467072 435134
rect 466400 434866 467072 434898
rect 493600 435454 494272 435486
rect 493600 435218 493658 435454
rect 493894 435218 493978 435454
rect 494214 435218 494272 435454
rect 493600 435134 494272 435218
rect 493600 434898 493658 435134
rect 493894 434898 493978 435134
rect 494214 434898 494272 435134
rect 493600 434866 494272 434898
rect 520800 435454 521472 435486
rect 520800 435218 520858 435454
rect 521094 435218 521178 435454
rect 521414 435218 521472 435454
rect 520800 435134 521472 435218
rect 520800 434898 520858 435134
rect 521094 434898 521178 435134
rect 521414 434898 521472 435134
rect 520800 434866 521472 434898
rect 548000 435454 548672 435486
rect 548000 435218 548058 435454
rect 548294 435218 548378 435454
rect 548614 435218 548672 435454
rect 548000 435134 548672 435218
rect 548000 434898 548058 435134
rect 548294 434898 548378 435134
rect 548614 434898 548672 435134
rect 548000 434866 548672 434898
rect 570260 435454 570880 435486
rect 570260 435218 570292 435454
rect 570528 435218 570612 435454
rect 570848 435218 570880 435454
rect 570260 435134 570880 435218
rect 570260 434898 570292 435134
rect 570528 434898 570612 435134
rect 570848 434898 570880 435134
rect 570260 434866 570880 434898
rect 7844 417454 8464 417486
rect 7844 417218 7876 417454
rect 8112 417218 8196 417454
rect 8432 417218 8464 417454
rect 7844 417134 8464 417218
rect 7844 416898 7876 417134
rect 8112 416898 8196 417134
rect 8432 416898 8464 417134
rect 7844 416866 8464 416898
rect 17600 417454 18272 417486
rect 17600 417218 17658 417454
rect 17894 417218 17978 417454
rect 18214 417218 18272 417454
rect 17600 417134 18272 417218
rect 17600 416898 17658 417134
rect 17894 416898 17978 417134
rect 18214 416898 18272 417134
rect 17600 416866 18272 416898
rect 44800 417454 45472 417486
rect 44800 417218 44858 417454
rect 45094 417218 45178 417454
rect 45414 417218 45472 417454
rect 44800 417134 45472 417218
rect 44800 416898 44858 417134
rect 45094 416898 45178 417134
rect 45414 416898 45472 417134
rect 44800 416866 45472 416898
rect 72000 417454 72672 417486
rect 72000 417218 72058 417454
rect 72294 417218 72378 417454
rect 72614 417218 72672 417454
rect 72000 417134 72672 417218
rect 72000 416898 72058 417134
rect 72294 416898 72378 417134
rect 72614 416898 72672 417134
rect 72000 416866 72672 416898
rect 99200 417454 99872 417486
rect 99200 417218 99258 417454
rect 99494 417218 99578 417454
rect 99814 417218 99872 417454
rect 99200 417134 99872 417218
rect 99200 416898 99258 417134
rect 99494 416898 99578 417134
rect 99814 416898 99872 417134
rect 99200 416866 99872 416898
rect 126400 417454 127072 417486
rect 126400 417218 126458 417454
rect 126694 417218 126778 417454
rect 127014 417218 127072 417454
rect 126400 417134 127072 417218
rect 126400 416898 126458 417134
rect 126694 416898 126778 417134
rect 127014 416898 127072 417134
rect 126400 416866 127072 416898
rect 153600 417454 154272 417486
rect 153600 417218 153658 417454
rect 153894 417218 153978 417454
rect 154214 417218 154272 417454
rect 153600 417134 154272 417218
rect 153600 416898 153658 417134
rect 153894 416898 153978 417134
rect 154214 416898 154272 417134
rect 153600 416866 154272 416898
rect 180800 417454 181472 417486
rect 180800 417218 180858 417454
rect 181094 417218 181178 417454
rect 181414 417218 181472 417454
rect 180800 417134 181472 417218
rect 180800 416898 180858 417134
rect 181094 416898 181178 417134
rect 181414 416898 181472 417134
rect 180800 416866 181472 416898
rect 208000 417454 208672 417486
rect 208000 417218 208058 417454
rect 208294 417218 208378 417454
rect 208614 417218 208672 417454
rect 208000 417134 208672 417218
rect 208000 416898 208058 417134
rect 208294 416898 208378 417134
rect 208614 416898 208672 417134
rect 208000 416866 208672 416898
rect 235200 417454 235872 417486
rect 235200 417218 235258 417454
rect 235494 417218 235578 417454
rect 235814 417218 235872 417454
rect 235200 417134 235872 417218
rect 235200 416898 235258 417134
rect 235494 416898 235578 417134
rect 235814 416898 235872 417134
rect 235200 416866 235872 416898
rect 262400 417454 263072 417486
rect 262400 417218 262458 417454
rect 262694 417218 262778 417454
rect 263014 417218 263072 417454
rect 262400 417134 263072 417218
rect 262400 416898 262458 417134
rect 262694 416898 262778 417134
rect 263014 416898 263072 417134
rect 262400 416866 263072 416898
rect 289600 417454 290272 417486
rect 289600 417218 289658 417454
rect 289894 417218 289978 417454
rect 290214 417218 290272 417454
rect 289600 417134 290272 417218
rect 289600 416898 289658 417134
rect 289894 416898 289978 417134
rect 290214 416898 290272 417134
rect 289600 416866 290272 416898
rect 316800 417454 317472 417486
rect 316800 417218 316858 417454
rect 317094 417218 317178 417454
rect 317414 417218 317472 417454
rect 316800 417134 317472 417218
rect 316800 416898 316858 417134
rect 317094 416898 317178 417134
rect 317414 416898 317472 417134
rect 316800 416866 317472 416898
rect 341763 417454 342123 417486
rect 341763 417218 341825 417454
rect 342061 417218 342123 417454
rect 341763 417134 342123 417218
rect 341763 416898 341825 417134
rect 342061 416898 342123 417134
rect 341763 416866 342123 416898
rect 440239 417454 440599 417486
rect 440239 417218 440301 417454
rect 440537 417218 440599 417454
rect 440239 417134 440599 417218
rect 440239 416898 440301 417134
rect 440537 416898 440599 417134
rect 440239 416866 440599 416898
rect 445735 417454 446095 417486
rect 445735 417218 445797 417454
rect 446033 417218 446095 417454
rect 445735 417134 446095 417218
rect 445735 416898 445797 417134
rect 446033 416898 446095 417134
rect 445735 416866 446095 416898
rect 544211 417454 544571 417486
rect 544211 417218 544273 417454
rect 544509 417218 544571 417454
rect 544211 417134 544571 417218
rect 544211 416898 544273 417134
rect 544509 416898 544571 417134
rect 544211 416866 544571 416898
rect 561600 417454 562272 417486
rect 561600 417218 561658 417454
rect 561894 417218 561978 417454
rect 562214 417218 562272 417454
rect 561600 417134 562272 417218
rect 561600 416898 561658 417134
rect 561894 416898 561978 417134
rect 562214 416898 562272 417134
rect 561600 416866 562272 416898
rect 571500 417454 572120 417486
rect 571500 417218 571532 417454
rect 571768 417218 571852 417454
rect 572088 417218 572120 417454
rect 571500 417134 572120 417218
rect 571500 416898 571532 417134
rect 571768 416898 571852 417134
rect 572088 416898 572120 417134
rect 571500 416866 572120 416898
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect 9084 399454 9704 399486
rect 9084 399218 9116 399454
rect 9352 399218 9436 399454
rect 9672 399218 9704 399454
rect 9084 399134 9704 399218
rect 9084 398898 9116 399134
rect 9352 398898 9436 399134
rect 9672 398898 9704 399134
rect 9084 398866 9704 398898
rect 31200 399454 31872 399486
rect 31200 399218 31258 399454
rect 31494 399218 31578 399454
rect 31814 399218 31872 399454
rect 31200 399134 31872 399218
rect 31200 398898 31258 399134
rect 31494 398898 31578 399134
rect 31814 398898 31872 399134
rect 31200 398866 31872 398898
rect 58400 399454 59072 399486
rect 58400 399218 58458 399454
rect 58694 399218 58778 399454
rect 59014 399218 59072 399454
rect 58400 399134 59072 399218
rect 58400 398898 58458 399134
rect 58694 398898 58778 399134
rect 59014 398898 59072 399134
rect 58400 398866 59072 398898
rect 85600 399454 86272 399486
rect 85600 399218 85658 399454
rect 85894 399218 85978 399454
rect 86214 399218 86272 399454
rect 85600 399134 86272 399218
rect 85600 398898 85658 399134
rect 85894 398898 85978 399134
rect 86214 398898 86272 399134
rect 85600 398866 86272 398898
rect 112800 399454 113472 399486
rect 112800 399218 112858 399454
rect 113094 399218 113178 399454
rect 113414 399218 113472 399454
rect 112800 399134 113472 399218
rect 112800 398898 112858 399134
rect 113094 398898 113178 399134
rect 113414 398898 113472 399134
rect 112800 398866 113472 398898
rect 140000 399454 140672 399486
rect 140000 399218 140058 399454
rect 140294 399218 140378 399454
rect 140614 399218 140672 399454
rect 140000 399134 140672 399218
rect 140000 398898 140058 399134
rect 140294 398898 140378 399134
rect 140614 398898 140672 399134
rect 140000 398866 140672 398898
rect 167200 399454 167872 399486
rect 167200 399218 167258 399454
rect 167494 399218 167578 399454
rect 167814 399218 167872 399454
rect 167200 399134 167872 399218
rect 167200 398898 167258 399134
rect 167494 398898 167578 399134
rect 167814 398898 167872 399134
rect 167200 398866 167872 398898
rect 194400 399454 195072 399486
rect 194400 399218 194458 399454
rect 194694 399218 194778 399454
rect 195014 399218 195072 399454
rect 194400 399134 195072 399218
rect 194400 398898 194458 399134
rect 194694 398898 194778 399134
rect 195014 398898 195072 399134
rect 194400 398866 195072 398898
rect 221600 399454 222272 399486
rect 221600 399218 221658 399454
rect 221894 399218 221978 399454
rect 222214 399218 222272 399454
rect 221600 399134 222272 399218
rect 221600 398898 221658 399134
rect 221894 398898 221978 399134
rect 222214 398898 222272 399134
rect 221600 398866 222272 398898
rect 248800 399454 249472 399486
rect 248800 399218 248858 399454
rect 249094 399218 249178 399454
rect 249414 399218 249472 399454
rect 248800 399134 249472 399218
rect 248800 398898 248858 399134
rect 249094 398898 249178 399134
rect 249414 398898 249472 399134
rect 248800 398866 249472 398898
rect 276000 399454 276672 399486
rect 276000 399218 276058 399454
rect 276294 399218 276378 399454
rect 276614 399218 276672 399454
rect 276000 399134 276672 399218
rect 276000 398898 276058 399134
rect 276294 398898 276378 399134
rect 276614 398898 276672 399134
rect 276000 398866 276672 398898
rect 303200 399454 303872 399486
rect 303200 399218 303258 399454
rect 303494 399218 303578 399454
rect 303814 399218 303872 399454
rect 303200 399134 303872 399218
rect 303200 398898 303258 399134
rect 303494 398898 303578 399134
rect 303814 398898 303872 399134
rect 303200 398866 303872 398898
rect 330400 399454 331072 399486
rect 330400 399218 330458 399454
rect 330694 399218 330778 399454
rect 331014 399218 331072 399454
rect 330400 399134 331072 399218
rect 330400 398898 330458 399134
rect 330694 398898 330778 399134
rect 331014 398898 331072 399134
rect 330400 398866 331072 398898
rect 342483 399454 342843 399486
rect 342483 399218 342545 399454
rect 342781 399218 342843 399454
rect 342483 399134 342843 399218
rect 342483 398898 342545 399134
rect 342781 398898 342843 399134
rect 342483 398866 342843 398898
rect 439519 399454 439879 399486
rect 439519 399218 439581 399454
rect 439817 399218 439879 399454
rect 439519 399134 439879 399218
rect 439519 398898 439581 399134
rect 439817 398898 439879 399134
rect 439519 398866 439879 398898
rect 446455 399454 446815 399486
rect 446455 399218 446517 399454
rect 446753 399218 446815 399454
rect 446455 399134 446815 399218
rect 446455 398898 446517 399134
rect 446753 398898 446815 399134
rect 446455 398866 446815 398898
rect 543491 399454 543851 399486
rect 543491 399218 543553 399454
rect 543789 399218 543851 399454
rect 543491 399134 543851 399218
rect 543491 398898 543553 399134
rect 543789 398898 543851 399134
rect 543491 398866 543851 398898
rect 548000 399454 548672 399486
rect 548000 399218 548058 399454
rect 548294 399218 548378 399454
rect 548614 399218 548672 399454
rect 548000 399134 548672 399218
rect 548000 398898 548058 399134
rect 548294 398898 548378 399134
rect 548614 398898 548672 399134
rect 548000 398866 548672 398898
rect 570260 399454 570880 399486
rect 570260 399218 570292 399454
rect 570528 399218 570612 399454
rect 570848 399218 570880 399454
rect 570260 399134 570880 399218
rect 570260 398898 570292 399134
rect 570528 398898 570612 399134
rect 570848 398898 570880 399134
rect 570260 398866 570880 398898
rect 7844 381454 8464 381486
rect 7844 381218 7876 381454
rect 8112 381218 8196 381454
rect 8432 381218 8464 381454
rect 7844 381134 8464 381218
rect 7844 380898 7876 381134
rect 8112 380898 8196 381134
rect 8432 380898 8464 381134
rect 7844 380866 8464 380898
rect 17600 381454 18272 381486
rect 17600 381218 17658 381454
rect 17894 381218 17978 381454
rect 18214 381218 18272 381454
rect 17600 381134 18272 381218
rect 17600 380898 17658 381134
rect 17894 380898 17978 381134
rect 18214 380898 18272 381134
rect 17600 380866 18272 380898
rect 44800 381454 45472 381486
rect 44800 381218 44858 381454
rect 45094 381218 45178 381454
rect 45414 381218 45472 381454
rect 44800 381134 45472 381218
rect 44800 380898 44858 381134
rect 45094 380898 45178 381134
rect 45414 380898 45472 381134
rect 44800 380866 45472 380898
rect 72000 381454 72672 381486
rect 72000 381218 72058 381454
rect 72294 381218 72378 381454
rect 72614 381218 72672 381454
rect 72000 381134 72672 381218
rect 72000 380898 72058 381134
rect 72294 380898 72378 381134
rect 72614 380898 72672 381134
rect 72000 380866 72672 380898
rect 99200 381454 99872 381486
rect 99200 381218 99258 381454
rect 99494 381218 99578 381454
rect 99814 381218 99872 381454
rect 99200 381134 99872 381218
rect 99200 380898 99258 381134
rect 99494 380898 99578 381134
rect 99814 380898 99872 381134
rect 99200 380866 99872 380898
rect 126400 381454 127072 381486
rect 126400 381218 126458 381454
rect 126694 381218 126778 381454
rect 127014 381218 127072 381454
rect 126400 381134 127072 381218
rect 126400 380898 126458 381134
rect 126694 380898 126778 381134
rect 127014 380898 127072 381134
rect 126400 380866 127072 380898
rect 153600 381454 154272 381486
rect 153600 381218 153658 381454
rect 153894 381218 153978 381454
rect 154214 381218 154272 381454
rect 153600 381134 154272 381218
rect 153600 380898 153658 381134
rect 153894 380898 153978 381134
rect 154214 380898 154272 381134
rect 153600 380866 154272 380898
rect 180800 381454 181472 381486
rect 180800 381218 180858 381454
rect 181094 381218 181178 381454
rect 181414 381218 181472 381454
rect 180800 381134 181472 381218
rect 180800 380898 180858 381134
rect 181094 380898 181178 381134
rect 181414 380898 181472 381134
rect 180800 380866 181472 380898
rect 208000 381454 208672 381486
rect 208000 381218 208058 381454
rect 208294 381218 208378 381454
rect 208614 381218 208672 381454
rect 208000 381134 208672 381218
rect 208000 380898 208058 381134
rect 208294 380898 208378 381134
rect 208614 380898 208672 381134
rect 208000 380866 208672 380898
rect 235200 381454 235872 381486
rect 235200 381218 235258 381454
rect 235494 381218 235578 381454
rect 235814 381218 235872 381454
rect 235200 381134 235872 381218
rect 235200 380898 235258 381134
rect 235494 380898 235578 381134
rect 235814 380898 235872 381134
rect 235200 380866 235872 380898
rect 262400 381454 263072 381486
rect 262400 381218 262458 381454
rect 262694 381218 262778 381454
rect 263014 381218 263072 381454
rect 262400 381134 263072 381218
rect 262400 380898 262458 381134
rect 262694 380898 262778 381134
rect 263014 380898 263072 381134
rect 262400 380866 263072 380898
rect 289600 381454 290272 381486
rect 289600 381218 289658 381454
rect 289894 381218 289978 381454
rect 290214 381218 290272 381454
rect 289600 381134 290272 381218
rect 289600 380898 289658 381134
rect 289894 380898 289978 381134
rect 290214 380898 290272 381134
rect 289600 380866 290272 380898
rect 316800 381454 317472 381486
rect 316800 381218 316858 381454
rect 317094 381218 317178 381454
rect 317414 381218 317472 381454
rect 316800 381134 317472 381218
rect 316800 380898 316858 381134
rect 317094 380898 317178 381134
rect 317414 380898 317472 381134
rect 316800 380866 317472 380898
rect 341763 381454 342123 381486
rect 341763 381218 341825 381454
rect 342061 381218 342123 381454
rect 341763 381134 342123 381218
rect 341763 380898 341825 381134
rect 342061 380898 342123 381134
rect 341763 380866 342123 380898
rect 440239 381454 440599 381486
rect 440239 381218 440301 381454
rect 440537 381218 440599 381454
rect 440239 381134 440599 381218
rect 440239 380898 440301 381134
rect 440537 380898 440599 381134
rect 440239 380866 440599 380898
rect 445735 381454 446095 381486
rect 445735 381218 445797 381454
rect 446033 381218 446095 381454
rect 445735 381134 446095 381218
rect 445735 380898 445797 381134
rect 446033 380898 446095 381134
rect 445735 380866 446095 380898
rect 544211 381454 544571 381486
rect 544211 381218 544273 381454
rect 544509 381218 544571 381454
rect 544211 381134 544571 381218
rect 544211 380898 544273 381134
rect 544509 380898 544571 381134
rect 544211 380866 544571 380898
rect 561600 381454 562272 381486
rect 561600 381218 561658 381454
rect 561894 381218 561978 381454
rect 562214 381218 562272 381454
rect 561600 381134 562272 381218
rect 561600 380898 561658 381134
rect 561894 380898 561978 381134
rect 562214 380898 562272 381134
rect 561600 380866 562272 380898
rect 571500 381454 572120 381486
rect 571500 381218 571532 381454
rect 571768 381218 571852 381454
rect 572088 381218 572120 381454
rect 571500 381134 572120 381218
rect 571500 380898 571532 381134
rect 571768 380898 571852 381134
rect 572088 380898 572120 381134
rect 571500 380866 572120 380898
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect 9084 363454 9704 363486
rect 9084 363218 9116 363454
rect 9352 363218 9436 363454
rect 9672 363218 9704 363454
rect 9084 363134 9704 363218
rect 9084 362898 9116 363134
rect 9352 362898 9436 363134
rect 9672 362898 9704 363134
rect 9084 362866 9704 362898
rect 31200 363454 31872 363486
rect 31200 363218 31258 363454
rect 31494 363218 31578 363454
rect 31814 363218 31872 363454
rect 31200 363134 31872 363218
rect 31200 362898 31258 363134
rect 31494 362898 31578 363134
rect 31814 362898 31872 363134
rect 31200 362866 31872 362898
rect 35555 363454 35915 363486
rect 35555 363218 35617 363454
rect 35853 363218 35915 363454
rect 35555 363134 35915 363218
rect 35555 362898 35617 363134
rect 35853 362898 35915 363134
rect 35555 362866 35915 362898
rect 132591 363454 132951 363486
rect 132591 363218 132653 363454
rect 132889 363218 132951 363454
rect 132591 363134 132951 363218
rect 132591 362898 132653 363134
rect 132889 362898 132951 363134
rect 132591 362866 132951 362898
rect 139527 363454 139887 363486
rect 139527 363218 139589 363454
rect 139825 363218 139887 363454
rect 139527 363134 139887 363218
rect 139527 362898 139589 363134
rect 139825 362898 139887 363134
rect 139527 362866 139887 362898
rect 236563 363454 236923 363486
rect 236563 363218 236625 363454
rect 236861 363218 236923 363454
rect 236563 363134 236923 363218
rect 236563 362898 236625 363134
rect 236861 362898 236923 363134
rect 236563 362866 236923 362898
rect 248800 363454 249472 363486
rect 248800 363218 248858 363454
rect 249094 363218 249178 363454
rect 249414 363218 249472 363454
rect 248800 363134 249472 363218
rect 248800 362898 248858 363134
rect 249094 362898 249178 363134
rect 249414 362898 249472 363134
rect 248800 362866 249472 362898
rect 276000 363454 276672 363486
rect 276000 363218 276058 363454
rect 276294 363218 276378 363454
rect 276614 363218 276672 363454
rect 276000 363134 276672 363218
rect 276000 362898 276058 363134
rect 276294 362898 276378 363134
rect 276614 362898 276672 363134
rect 276000 362866 276672 362898
rect 303200 363454 303872 363486
rect 303200 363218 303258 363454
rect 303494 363218 303578 363454
rect 303814 363218 303872 363454
rect 303200 363134 303872 363218
rect 303200 362898 303258 363134
rect 303494 362898 303578 363134
rect 303814 362898 303872 363134
rect 303200 362866 303872 362898
rect 330400 363454 331072 363486
rect 330400 363218 330458 363454
rect 330694 363218 330778 363454
rect 331014 363218 331072 363454
rect 330400 363134 331072 363218
rect 330400 362898 330458 363134
rect 330694 362898 330778 363134
rect 331014 362898 331072 363134
rect 330400 362866 331072 362898
rect 342483 363454 342843 363486
rect 342483 363218 342545 363454
rect 342781 363218 342843 363454
rect 342483 363134 342843 363218
rect 342483 362898 342545 363134
rect 342781 362898 342843 363134
rect 342483 362866 342843 362898
rect 439519 363454 439879 363486
rect 439519 363218 439581 363454
rect 439817 363218 439879 363454
rect 439519 363134 439879 363218
rect 439519 362898 439581 363134
rect 439817 362898 439879 363134
rect 439519 362866 439879 362898
rect 446455 363454 446815 363486
rect 446455 363218 446517 363454
rect 446753 363218 446815 363454
rect 446455 363134 446815 363218
rect 446455 362898 446517 363134
rect 446753 362898 446815 363134
rect 446455 362866 446815 362898
rect 543491 363454 543851 363486
rect 543491 363218 543553 363454
rect 543789 363218 543851 363454
rect 543491 363134 543851 363218
rect 543491 362898 543553 363134
rect 543789 362898 543851 363134
rect 543491 362866 543851 362898
rect 548000 363454 548672 363486
rect 548000 363218 548058 363454
rect 548294 363218 548378 363454
rect 548614 363218 548672 363454
rect 548000 363134 548672 363218
rect 548000 362898 548058 363134
rect 548294 362898 548378 363134
rect 548614 362898 548672 363134
rect 548000 362866 548672 362898
rect 570260 363454 570880 363486
rect 570260 363218 570292 363454
rect 570528 363218 570612 363454
rect 570848 363218 570880 363454
rect 570260 363134 570880 363218
rect 570260 362898 570292 363134
rect 570528 362898 570612 363134
rect 570848 362898 570880 363134
rect 570260 362866 570880 362898
rect 7844 345454 8464 345486
rect 7844 345218 7876 345454
rect 8112 345218 8196 345454
rect 8432 345218 8464 345454
rect 7844 345134 8464 345218
rect 7844 344898 7876 345134
rect 8112 344898 8196 345134
rect 8432 344898 8464 345134
rect 7844 344866 8464 344898
rect 17600 345454 18272 345486
rect 17600 345218 17658 345454
rect 17894 345218 17978 345454
rect 18214 345218 18272 345454
rect 17600 345134 18272 345218
rect 17600 344898 17658 345134
rect 17894 344898 17978 345134
rect 18214 344898 18272 345134
rect 17600 344866 18272 344898
rect 34835 345454 35195 345486
rect 34835 345218 34897 345454
rect 35133 345218 35195 345454
rect 34835 345134 35195 345218
rect 34835 344898 34897 345134
rect 35133 344898 35195 345134
rect 34835 344866 35195 344898
rect 133311 345454 133671 345486
rect 133311 345218 133373 345454
rect 133609 345218 133671 345454
rect 133311 345134 133671 345218
rect 133311 344898 133373 345134
rect 133609 344898 133671 345134
rect 133311 344866 133671 344898
rect 138807 345454 139167 345486
rect 138807 345218 138869 345454
rect 139105 345218 139167 345454
rect 138807 345134 139167 345218
rect 138807 344898 138869 345134
rect 139105 344898 139167 345134
rect 138807 344866 139167 344898
rect 237283 345454 237643 345486
rect 237283 345218 237345 345454
rect 237581 345218 237643 345454
rect 237283 345134 237643 345218
rect 237283 344898 237345 345134
rect 237581 344898 237643 345134
rect 237283 344866 237643 344898
rect 262400 345454 263072 345486
rect 262400 345218 262458 345454
rect 262694 345218 262778 345454
rect 263014 345218 263072 345454
rect 262400 345134 263072 345218
rect 262400 344898 262458 345134
rect 262694 344898 262778 345134
rect 263014 344898 263072 345134
rect 262400 344866 263072 344898
rect 289600 345454 290272 345486
rect 289600 345218 289658 345454
rect 289894 345218 289978 345454
rect 290214 345218 290272 345454
rect 289600 345134 290272 345218
rect 289600 344898 289658 345134
rect 289894 344898 289978 345134
rect 290214 344898 290272 345134
rect 289600 344866 290272 344898
rect 316800 345454 317472 345486
rect 316800 345218 316858 345454
rect 317094 345218 317178 345454
rect 317414 345218 317472 345454
rect 316800 345134 317472 345218
rect 316800 344898 316858 345134
rect 317094 344898 317178 345134
rect 317414 344898 317472 345134
rect 316800 344866 317472 344898
rect 341763 345454 342123 345486
rect 341763 345218 341825 345454
rect 342061 345218 342123 345454
rect 341763 345134 342123 345218
rect 341763 344898 341825 345134
rect 342061 344898 342123 345134
rect 341763 344866 342123 344898
rect 440239 345454 440599 345486
rect 440239 345218 440301 345454
rect 440537 345218 440599 345454
rect 440239 345134 440599 345218
rect 440239 344898 440301 345134
rect 440537 344898 440599 345134
rect 440239 344866 440599 344898
rect 445735 345454 446095 345486
rect 445735 345218 445797 345454
rect 446033 345218 446095 345454
rect 445735 345134 446095 345218
rect 445735 344898 445797 345134
rect 446033 344898 446095 345134
rect 445735 344866 446095 344898
rect 544211 345454 544571 345486
rect 544211 345218 544273 345454
rect 544509 345218 544571 345454
rect 544211 345134 544571 345218
rect 544211 344898 544273 345134
rect 544509 344898 544571 345134
rect 544211 344866 544571 344898
rect 561600 345454 562272 345486
rect 561600 345218 561658 345454
rect 561894 345218 561978 345454
rect 562214 345218 562272 345454
rect 561600 345134 562272 345218
rect 561600 344898 561658 345134
rect 561894 344898 561978 345134
rect 562214 344898 562272 345134
rect 561600 344866 562272 344898
rect 571500 345454 572120 345486
rect 571500 345218 571532 345454
rect 571768 345218 571852 345454
rect 572088 345218 572120 345454
rect 571500 345134 572120 345218
rect 571500 344898 571532 345134
rect 571768 344898 571852 345134
rect 572088 344898 572120 345134
rect 571500 344866 572120 344898
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect 9084 327454 9704 327486
rect 9084 327218 9116 327454
rect 9352 327218 9436 327454
rect 9672 327218 9704 327454
rect 9084 327134 9704 327218
rect 9084 326898 9116 327134
rect 9352 326898 9436 327134
rect 9672 326898 9704 327134
rect 9084 326866 9704 326898
rect 31200 327454 31872 327486
rect 31200 327218 31258 327454
rect 31494 327218 31578 327454
rect 31814 327218 31872 327454
rect 31200 327134 31872 327218
rect 31200 326898 31258 327134
rect 31494 326898 31578 327134
rect 31814 326898 31872 327134
rect 31200 326866 31872 326898
rect 35555 327454 35915 327486
rect 35555 327218 35617 327454
rect 35853 327218 35915 327454
rect 35555 327134 35915 327218
rect 35555 326898 35617 327134
rect 35853 326898 35915 327134
rect 35555 326866 35915 326898
rect 132591 327454 132951 327486
rect 132591 327218 132653 327454
rect 132889 327218 132951 327454
rect 132591 327134 132951 327218
rect 132591 326898 132653 327134
rect 132889 326898 132951 327134
rect 132591 326866 132951 326898
rect 139527 327454 139887 327486
rect 139527 327218 139589 327454
rect 139825 327218 139887 327454
rect 139527 327134 139887 327218
rect 139527 326898 139589 327134
rect 139825 326898 139887 327134
rect 139527 326866 139887 326898
rect 236563 327454 236923 327486
rect 236563 327218 236625 327454
rect 236861 327218 236923 327454
rect 236563 327134 236923 327218
rect 236563 326898 236625 327134
rect 236861 326898 236923 327134
rect 236563 326866 236923 326898
rect 248800 327454 249472 327486
rect 248800 327218 248858 327454
rect 249094 327218 249178 327454
rect 249414 327218 249472 327454
rect 248800 327134 249472 327218
rect 248800 326898 248858 327134
rect 249094 326898 249178 327134
rect 249414 326898 249472 327134
rect 248800 326866 249472 326898
rect 276000 327454 276672 327486
rect 276000 327218 276058 327454
rect 276294 327218 276378 327454
rect 276614 327218 276672 327454
rect 276000 327134 276672 327218
rect 276000 326898 276058 327134
rect 276294 326898 276378 327134
rect 276614 326898 276672 327134
rect 276000 326866 276672 326898
rect 303200 327454 303872 327486
rect 303200 327218 303258 327454
rect 303494 327218 303578 327454
rect 303814 327218 303872 327454
rect 303200 327134 303872 327218
rect 303200 326898 303258 327134
rect 303494 326898 303578 327134
rect 303814 326898 303872 327134
rect 303200 326866 303872 326898
rect 330400 327454 331072 327486
rect 330400 327218 330458 327454
rect 330694 327218 330778 327454
rect 331014 327218 331072 327454
rect 330400 327134 331072 327218
rect 330400 326898 330458 327134
rect 330694 326898 330778 327134
rect 331014 326898 331072 327134
rect 330400 326866 331072 326898
rect 342483 327454 342843 327486
rect 342483 327218 342545 327454
rect 342781 327218 342843 327454
rect 342483 327134 342843 327218
rect 342483 326898 342545 327134
rect 342781 326898 342843 327134
rect 342483 326866 342843 326898
rect 446455 327454 446815 327486
rect 446455 327218 446517 327454
rect 446753 327218 446815 327454
rect 446455 327134 446815 327218
rect 446455 326898 446517 327134
rect 446753 326898 446815 327134
rect 446455 326866 446815 326898
rect 543491 327454 543851 327486
rect 543491 327218 543553 327454
rect 543789 327218 543851 327454
rect 543491 327134 543851 327218
rect 543491 326898 543553 327134
rect 543789 326898 543851 327134
rect 543491 326866 543851 326898
rect 548000 327454 548672 327486
rect 548000 327218 548058 327454
rect 548294 327218 548378 327454
rect 548614 327218 548672 327454
rect 548000 327134 548672 327218
rect 548000 326898 548058 327134
rect 548294 326898 548378 327134
rect 548614 326898 548672 327134
rect 548000 326866 548672 326898
rect 570260 327454 570880 327486
rect 570260 327218 570292 327454
rect 570528 327218 570612 327454
rect 570848 327218 570880 327454
rect 570260 327134 570880 327218
rect 570260 326898 570292 327134
rect 570528 326898 570612 327134
rect 570848 326898 570880 327134
rect 570260 326866 570880 326898
rect 7844 309454 8464 309486
rect 7844 309218 7876 309454
rect 8112 309218 8196 309454
rect 8432 309218 8464 309454
rect 7844 309134 8464 309218
rect 7844 308898 7876 309134
rect 8112 308898 8196 309134
rect 8432 308898 8464 309134
rect 7844 308866 8464 308898
rect 17600 309454 18272 309486
rect 17600 309218 17658 309454
rect 17894 309218 17978 309454
rect 18214 309218 18272 309454
rect 17600 309134 18272 309218
rect 17600 308898 17658 309134
rect 17894 308898 17978 309134
rect 18214 308898 18272 309134
rect 17600 308866 18272 308898
rect 34835 309454 35195 309486
rect 34835 309218 34897 309454
rect 35133 309218 35195 309454
rect 34835 309134 35195 309218
rect 34835 308898 34897 309134
rect 35133 308898 35195 309134
rect 34835 308866 35195 308898
rect 133311 309454 133671 309486
rect 133311 309218 133373 309454
rect 133609 309218 133671 309454
rect 133311 309134 133671 309218
rect 133311 308898 133373 309134
rect 133609 308898 133671 309134
rect 133311 308866 133671 308898
rect 138807 309454 139167 309486
rect 138807 309218 138869 309454
rect 139105 309218 139167 309454
rect 138807 309134 139167 309218
rect 138807 308898 138869 309134
rect 139105 308898 139167 309134
rect 138807 308866 139167 308898
rect 237283 309454 237643 309486
rect 237283 309218 237345 309454
rect 237581 309218 237643 309454
rect 237283 309134 237643 309218
rect 237283 308898 237345 309134
rect 237581 308898 237643 309134
rect 237283 308866 237643 308898
rect 262400 309454 263072 309486
rect 262400 309218 262458 309454
rect 262694 309218 262778 309454
rect 263014 309218 263072 309454
rect 262400 309134 263072 309218
rect 262400 308898 262458 309134
rect 262694 308898 262778 309134
rect 263014 308898 263072 309134
rect 262400 308866 263072 308898
rect 289600 309454 290272 309486
rect 289600 309218 289658 309454
rect 289894 309218 289978 309454
rect 290214 309218 290272 309454
rect 289600 309134 290272 309218
rect 289600 308898 289658 309134
rect 289894 308898 289978 309134
rect 290214 308898 290272 309134
rect 289600 308866 290272 308898
rect 316800 309454 317472 309486
rect 316800 309218 316858 309454
rect 317094 309218 317178 309454
rect 317414 309218 317472 309454
rect 316800 309134 317472 309218
rect 316800 308898 316858 309134
rect 317094 308898 317178 309134
rect 317414 308898 317472 309134
rect 316800 308866 317472 308898
rect 341763 309454 342123 309486
rect 341763 309218 341825 309454
rect 342061 309218 342123 309454
rect 341763 309134 342123 309218
rect 341763 308898 341825 309134
rect 342061 308898 342123 309134
rect 341763 308866 342123 308898
rect 440239 309454 440599 309486
rect 440239 309218 440301 309454
rect 440537 309218 440599 309454
rect 440239 309134 440599 309218
rect 440239 308898 440301 309134
rect 440537 308898 440599 309134
rect 440239 308866 440599 308898
rect 445735 309454 446095 309486
rect 445735 309218 445797 309454
rect 446033 309218 446095 309454
rect 445735 309134 446095 309218
rect 445735 308898 445797 309134
rect 446033 308898 446095 309134
rect 445735 308866 446095 308898
rect 544211 309454 544571 309486
rect 544211 309218 544273 309454
rect 544509 309218 544571 309454
rect 544211 309134 544571 309218
rect 544211 308898 544273 309134
rect 544509 308898 544571 309134
rect 544211 308866 544571 308898
rect 561600 309454 562272 309486
rect 561600 309218 561658 309454
rect 561894 309218 561978 309454
rect 562214 309218 562272 309454
rect 561600 309134 562272 309218
rect 561600 308898 561658 309134
rect 561894 308898 561978 309134
rect 562214 308898 562272 309134
rect 561600 308866 562272 308898
rect 571500 309454 572120 309486
rect 571500 309218 571532 309454
rect 571768 309218 571852 309454
rect 572088 309218 572120 309454
rect 571500 309134 572120 309218
rect 571500 308898 571532 309134
rect 571768 308898 571852 309134
rect 572088 308898 572120 309134
rect 571500 308866 572120 308898
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect 9084 291454 9704 291486
rect 9084 291218 9116 291454
rect 9352 291218 9436 291454
rect 9672 291218 9704 291454
rect 9084 291134 9704 291218
rect 9084 290898 9116 291134
rect 9352 290898 9436 291134
rect 9672 290898 9704 291134
rect 9084 290866 9704 290898
rect 31200 291454 31872 291486
rect 31200 291218 31258 291454
rect 31494 291218 31578 291454
rect 31814 291218 31872 291454
rect 31200 291134 31872 291218
rect 31200 290898 31258 291134
rect 31494 290898 31578 291134
rect 31814 290898 31872 291134
rect 31200 290866 31872 290898
rect 35555 291454 35915 291486
rect 35555 291218 35617 291454
rect 35853 291218 35915 291454
rect 35555 291134 35915 291218
rect 35555 290898 35617 291134
rect 35853 290898 35915 291134
rect 35555 290866 35915 290898
rect 132591 291454 132951 291486
rect 132591 291218 132653 291454
rect 132889 291218 132951 291454
rect 132591 291134 132951 291218
rect 132591 290898 132653 291134
rect 132889 290898 132951 291134
rect 132591 290866 132951 290898
rect 139527 291454 139887 291486
rect 139527 291218 139589 291454
rect 139825 291218 139887 291454
rect 139527 291134 139887 291218
rect 139527 290898 139589 291134
rect 139825 290898 139887 291134
rect 139527 290866 139887 290898
rect 236563 291454 236923 291486
rect 236563 291218 236625 291454
rect 236861 291218 236923 291454
rect 236563 291134 236923 291218
rect 236563 290898 236625 291134
rect 236861 290898 236923 291134
rect 236563 290866 236923 290898
rect 248800 291454 249472 291486
rect 248800 291218 248858 291454
rect 249094 291218 249178 291454
rect 249414 291218 249472 291454
rect 248800 291134 249472 291218
rect 248800 290898 248858 291134
rect 249094 290898 249178 291134
rect 249414 290898 249472 291134
rect 248800 290866 249472 290898
rect 276000 291454 276672 291486
rect 276000 291218 276058 291454
rect 276294 291218 276378 291454
rect 276614 291218 276672 291454
rect 276000 291134 276672 291218
rect 276000 290898 276058 291134
rect 276294 290898 276378 291134
rect 276614 290898 276672 291134
rect 276000 290866 276672 290898
rect 303200 291454 303872 291486
rect 303200 291218 303258 291454
rect 303494 291218 303578 291454
rect 303814 291218 303872 291454
rect 303200 291134 303872 291218
rect 303200 290898 303258 291134
rect 303494 290898 303578 291134
rect 303814 290898 303872 291134
rect 303200 290866 303872 290898
rect 330400 291454 331072 291486
rect 330400 291218 330458 291454
rect 330694 291218 330778 291454
rect 331014 291218 331072 291454
rect 330400 291134 331072 291218
rect 330400 290898 330458 291134
rect 330694 290898 330778 291134
rect 331014 290898 331072 291134
rect 330400 290866 331072 290898
rect 342483 291454 342843 291486
rect 342483 291218 342545 291454
rect 342781 291218 342843 291454
rect 342483 291134 342843 291218
rect 342483 290898 342545 291134
rect 342781 290898 342843 291134
rect 342483 290866 342843 290898
rect 439519 291454 439879 291486
rect 439519 291218 439581 291454
rect 439817 291218 439879 291454
rect 439519 291134 439879 291218
rect 439519 290898 439581 291134
rect 439817 290898 439879 291134
rect 439519 290866 439879 290898
rect 446455 291454 446815 291486
rect 446455 291218 446517 291454
rect 446753 291218 446815 291454
rect 446455 291134 446815 291218
rect 446455 290898 446517 291134
rect 446753 290898 446815 291134
rect 446455 290866 446815 290898
rect 543491 291454 543851 291486
rect 543491 291218 543553 291454
rect 543789 291218 543851 291454
rect 543491 291134 543851 291218
rect 543491 290898 543553 291134
rect 543789 290898 543851 291134
rect 543491 290866 543851 290898
rect 548000 291454 548672 291486
rect 548000 291218 548058 291454
rect 548294 291218 548378 291454
rect 548614 291218 548672 291454
rect 548000 291134 548672 291218
rect 548000 290898 548058 291134
rect 548294 290898 548378 291134
rect 548614 290898 548672 291134
rect 548000 290866 548672 290898
rect 570260 291454 570880 291486
rect 570260 291218 570292 291454
rect 570528 291218 570612 291454
rect 570848 291218 570880 291454
rect 570260 291134 570880 291218
rect 570260 290898 570292 291134
rect 570528 290898 570612 291134
rect 570848 290898 570880 291134
rect 570260 290866 570880 290898
rect 7844 273454 8464 273486
rect 7844 273218 7876 273454
rect 8112 273218 8196 273454
rect 8432 273218 8464 273454
rect 7844 273134 8464 273218
rect 7844 272898 7876 273134
rect 8112 272898 8196 273134
rect 8432 272898 8464 273134
rect 7844 272866 8464 272898
rect 17600 273454 18272 273486
rect 17600 273218 17658 273454
rect 17894 273218 17978 273454
rect 18214 273218 18272 273454
rect 17600 273134 18272 273218
rect 17600 272898 17658 273134
rect 17894 272898 17978 273134
rect 18214 272898 18272 273134
rect 17600 272866 18272 272898
rect 44800 273454 45472 273486
rect 44800 273218 44858 273454
rect 45094 273218 45178 273454
rect 45414 273218 45472 273454
rect 44800 273134 45472 273218
rect 44800 272898 44858 273134
rect 45094 272898 45178 273134
rect 45414 272898 45472 273134
rect 44800 272866 45472 272898
rect 72000 273454 72672 273486
rect 72000 273218 72058 273454
rect 72294 273218 72378 273454
rect 72614 273218 72672 273454
rect 72000 273134 72672 273218
rect 72000 272898 72058 273134
rect 72294 272898 72378 273134
rect 72614 272898 72672 273134
rect 72000 272866 72672 272898
rect 99200 273454 99872 273486
rect 99200 273218 99258 273454
rect 99494 273218 99578 273454
rect 99814 273218 99872 273454
rect 99200 273134 99872 273218
rect 99200 272898 99258 273134
rect 99494 272898 99578 273134
rect 99814 272898 99872 273134
rect 99200 272866 99872 272898
rect 126400 273454 127072 273486
rect 126400 273218 126458 273454
rect 126694 273218 126778 273454
rect 127014 273218 127072 273454
rect 126400 273134 127072 273218
rect 126400 272898 126458 273134
rect 126694 272898 126778 273134
rect 127014 272898 127072 273134
rect 126400 272866 127072 272898
rect 153600 273454 154272 273486
rect 153600 273218 153658 273454
rect 153894 273218 153978 273454
rect 154214 273218 154272 273454
rect 153600 273134 154272 273218
rect 153600 272898 153658 273134
rect 153894 272898 153978 273134
rect 154214 272898 154272 273134
rect 153600 272866 154272 272898
rect 180800 273454 181472 273486
rect 180800 273218 180858 273454
rect 181094 273218 181178 273454
rect 181414 273218 181472 273454
rect 180800 273134 181472 273218
rect 180800 272898 180858 273134
rect 181094 272898 181178 273134
rect 181414 272898 181472 273134
rect 180800 272866 181472 272898
rect 208000 273454 208672 273486
rect 208000 273218 208058 273454
rect 208294 273218 208378 273454
rect 208614 273218 208672 273454
rect 208000 273134 208672 273218
rect 208000 272898 208058 273134
rect 208294 272898 208378 273134
rect 208614 272898 208672 273134
rect 208000 272866 208672 272898
rect 235200 273454 235872 273486
rect 235200 273218 235258 273454
rect 235494 273218 235578 273454
rect 235814 273218 235872 273454
rect 235200 273134 235872 273218
rect 235200 272898 235258 273134
rect 235494 272898 235578 273134
rect 235814 272898 235872 273134
rect 235200 272866 235872 272898
rect 262400 273454 263072 273486
rect 262400 273218 262458 273454
rect 262694 273218 262778 273454
rect 263014 273218 263072 273454
rect 262400 273134 263072 273218
rect 262400 272898 262458 273134
rect 262694 272898 262778 273134
rect 263014 272898 263072 273134
rect 262400 272866 263072 272898
rect 289600 273454 290272 273486
rect 289600 273218 289658 273454
rect 289894 273218 289978 273454
rect 290214 273218 290272 273454
rect 289600 273134 290272 273218
rect 289600 272898 289658 273134
rect 289894 272898 289978 273134
rect 290214 272898 290272 273134
rect 289600 272866 290272 272898
rect 316800 273454 317472 273486
rect 316800 273218 316858 273454
rect 317094 273218 317178 273454
rect 317414 273218 317472 273454
rect 316800 273134 317472 273218
rect 316800 272898 316858 273134
rect 317094 272898 317178 273134
rect 317414 272898 317472 273134
rect 316800 272866 317472 272898
rect 341763 273454 342123 273486
rect 341763 273218 341825 273454
rect 342061 273218 342123 273454
rect 341763 273134 342123 273218
rect 341763 272898 341825 273134
rect 342061 272898 342123 273134
rect 341763 272866 342123 272898
rect 440239 273454 440599 273486
rect 440239 273218 440301 273454
rect 440537 273218 440599 273454
rect 440239 273134 440599 273218
rect 440239 272898 440301 273134
rect 440537 272898 440599 273134
rect 440239 272866 440599 272898
rect 445735 273454 446095 273486
rect 445735 273218 445797 273454
rect 446033 273218 446095 273454
rect 445735 273134 446095 273218
rect 445735 272898 445797 273134
rect 446033 272898 446095 273134
rect 445735 272866 446095 272898
rect 544211 273454 544571 273486
rect 544211 273218 544273 273454
rect 544509 273218 544571 273454
rect 544211 273134 544571 273218
rect 544211 272898 544273 273134
rect 544509 272898 544571 273134
rect 544211 272866 544571 272898
rect 561600 273454 562272 273486
rect 561600 273218 561658 273454
rect 561894 273218 561978 273454
rect 562214 273218 562272 273454
rect 561600 273134 562272 273218
rect 561600 272898 561658 273134
rect 561894 272898 561978 273134
rect 562214 272898 562272 273134
rect 561600 272866 562272 272898
rect 571500 273454 572120 273486
rect 571500 273218 571532 273454
rect 571768 273218 571852 273454
rect 572088 273218 572120 273454
rect 571500 273134 572120 273218
rect 571500 272898 571532 273134
rect 571768 272898 571852 273134
rect 572088 272898 572120 273134
rect 571500 272866 572120 272898
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect 9084 255454 9704 255486
rect 9084 255218 9116 255454
rect 9352 255218 9436 255454
rect 9672 255218 9704 255454
rect 9084 255134 9704 255218
rect 9084 254898 9116 255134
rect 9352 254898 9436 255134
rect 9672 254898 9704 255134
rect 9084 254866 9704 254898
rect 31200 255454 31872 255486
rect 31200 255218 31258 255454
rect 31494 255218 31578 255454
rect 31814 255218 31872 255454
rect 31200 255134 31872 255218
rect 31200 254898 31258 255134
rect 31494 254898 31578 255134
rect 31814 254898 31872 255134
rect 31200 254866 31872 254898
rect 58400 255454 59072 255486
rect 58400 255218 58458 255454
rect 58694 255218 58778 255454
rect 59014 255218 59072 255454
rect 58400 255134 59072 255218
rect 58400 254898 58458 255134
rect 58694 254898 58778 255134
rect 59014 254898 59072 255134
rect 58400 254866 59072 254898
rect 85600 255454 86272 255486
rect 85600 255218 85658 255454
rect 85894 255218 85978 255454
rect 86214 255218 86272 255454
rect 85600 255134 86272 255218
rect 85600 254898 85658 255134
rect 85894 254898 85978 255134
rect 86214 254898 86272 255134
rect 85600 254866 86272 254898
rect 112800 255454 113472 255486
rect 112800 255218 112858 255454
rect 113094 255218 113178 255454
rect 113414 255218 113472 255454
rect 112800 255134 113472 255218
rect 112800 254898 112858 255134
rect 113094 254898 113178 255134
rect 113414 254898 113472 255134
rect 112800 254866 113472 254898
rect 140000 255454 140672 255486
rect 140000 255218 140058 255454
rect 140294 255218 140378 255454
rect 140614 255218 140672 255454
rect 140000 255134 140672 255218
rect 140000 254898 140058 255134
rect 140294 254898 140378 255134
rect 140614 254898 140672 255134
rect 140000 254866 140672 254898
rect 167200 255454 167872 255486
rect 167200 255218 167258 255454
rect 167494 255218 167578 255454
rect 167814 255218 167872 255454
rect 167200 255134 167872 255218
rect 167200 254898 167258 255134
rect 167494 254898 167578 255134
rect 167814 254898 167872 255134
rect 167200 254866 167872 254898
rect 194400 255454 195072 255486
rect 194400 255218 194458 255454
rect 194694 255218 194778 255454
rect 195014 255218 195072 255454
rect 194400 255134 195072 255218
rect 194400 254898 194458 255134
rect 194694 254898 194778 255134
rect 195014 254898 195072 255134
rect 194400 254866 195072 254898
rect 221600 255454 222272 255486
rect 221600 255218 221658 255454
rect 221894 255218 221978 255454
rect 222214 255218 222272 255454
rect 221600 255134 222272 255218
rect 221600 254898 221658 255134
rect 221894 254898 221978 255134
rect 222214 254898 222272 255134
rect 221600 254866 222272 254898
rect 248800 255454 249472 255486
rect 248800 255218 248858 255454
rect 249094 255218 249178 255454
rect 249414 255218 249472 255454
rect 248800 255134 249472 255218
rect 248800 254898 248858 255134
rect 249094 254898 249178 255134
rect 249414 254898 249472 255134
rect 248800 254866 249472 254898
rect 276000 255454 276672 255486
rect 276000 255218 276058 255454
rect 276294 255218 276378 255454
rect 276614 255218 276672 255454
rect 276000 255134 276672 255218
rect 276000 254898 276058 255134
rect 276294 254898 276378 255134
rect 276614 254898 276672 255134
rect 276000 254866 276672 254898
rect 303200 255454 303872 255486
rect 303200 255218 303258 255454
rect 303494 255218 303578 255454
rect 303814 255218 303872 255454
rect 303200 255134 303872 255218
rect 303200 254898 303258 255134
rect 303494 254898 303578 255134
rect 303814 254898 303872 255134
rect 303200 254866 303872 254898
rect 330400 255454 331072 255486
rect 330400 255218 330458 255454
rect 330694 255218 330778 255454
rect 331014 255218 331072 255454
rect 330400 255134 331072 255218
rect 330400 254898 330458 255134
rect 330694 254898 330778 255134
rect 331014 254898 331072 255134
rect 330400 254866 331072 254898
rect 342483 255454 342843 255486
rect 342483 255218 342545 255454
rect 342781 255218 342843 255454
rect 342483 255134 342843 255218
rect 342483 254898 342545 255134
rect 342781 254898 342843 255134
rect 342483 254866 342843 254898
rect 439519 255454 439879 255486
rect 439519 255218 439581 255454
rect 439817 255218 439879 255454
rect 439519 255134 439879 255218
rect 439519 254898 439581 255134
rect 439817 254898 439879 255134
rect 439519 254866 439879 254898
rect 446455 255454 446815 255486
rect 446455 255218 446517 255454
rect 446753 255218 446815 255454
rect 446455 255134 446815 255218
rect 446455 254898 446517 255134
rect 446753 254898 446815 255134
rect 446455 254866 446815 254898
rect 543491 255454 543851 255486
rect 543491 255218 543553 255454
rect 543789 255218 543851 255454
rect 543491 255134 543851 255218
rect 543491 254898 543553 255134
rect 543789 254898 543851 255134
rect 543491 254866 543851 254898
rect 548000 255454 548672 255486
rect 548000 255218 548058 255454
rect 548294 255218 548378 255454
rect 548614 255218 548672 255454
rect 548000 255134 548672 255218
rect 548000 254898 548058 255134
rect 548294 254898 548378 255134
rect 548614 254898 548672 255134
rect 548000 254866 548672 254898
rect 570260 255454 570880 255486
rect 570260 255218 570292 255454
rect 570528 255218 570612 255454
rect 570848 255218 570880 255454
rect 570260 255134 570880 255218
rect 570260 254898 570292 255134
rect 570528 254898 570612 255134
rect 570848 254898 570880 255134
rect 570260 254866 570880 254898
rect 7844 237454 8464 237486
rect 7844 237218 7876 237454
rect 8112 237218 8196 237454
rect 8432 237218 8464 237454
rect 7844 237134 8464 237218
rect 7844 236898 7876 237134
rect 8112 236898 8196 237134
rect 8432 236898 8464 237134
rect 7844 236866 8464 236898
rect 17600 237454 18272 237486
rect 17600 237218 17658 237454
rect 17894 237218 17978 237454
rect 18214 237218 18272 237454
rect 17600 237134 18272 237218
rect 17600 236898 17658 237134
rect 17894 236898 17978 237134
rect 18214 236898 18272 237134
rect 17600 236866 18272 236898
rect 44800 237454 45472 237486
rect 44800 237218 44858 237454
rect 45094 237218 45178 237454
rect 45414 237218 45472 237454
rect 44800 237134 45472 237218
rect 44800 236898 44858 237134
rect 45094 236898 45178 237134
rect 45414 236898 45472 237134
rect 44800 236866 45472 236898
rect 72000 237454 72672 237486
rect 72000 237218 72058 237454
rect 72294 237218 72378 237454
rect 72614 237218 72672 237454
rect 72000 237134 72672 237218
rect 72000 236898 72058 237134
rect 72294 236898 72378 237134
rect 72614 236898 72672 237134
rect 72000 236866 72672 236898
rect 99200 237454 99872 237486
rect 99200 237218 99258 237454
rect 99494 237218 99578 237454
rect 99814 237218 99872 237454
rect 99200 237134 99872 237218
rect 99200 236898 99258 237134
rect 99494 236898 99578 237134
rect 99814 236898 99872 237134
rect 99200 236866 99872 236898
rect 126400 237454 127072 237486
rect 126400 237218 126458 237454
rect 126694 237218 126778 237454
rect 127014 237218 127072 237454
rect 126400 237134 127072 237218
rect 126400 236898 126458 237134
rect 126694 236898 126778 237134
rect 127014 236898 127072 237134
rect 126400 236866 127072 236898
rect 153600 237454 154272 237486
rect 153600 237218 153658 237454
rect 153894 237218 153978 237454
rect 154214 237218 154272 237454
rect 153600 237134 154272 237218
rect 153600 236898 153658 237134
rect 153894 236898 153978 237134
rect 154214 236898 154272 237134
rect 153600 236866 154272 236898
rect 180800 237454 181472 237486
rect 180800 237218 180858 237454
rect 181094 237218 181178 237454
rect 181414 237218 181472 237454
rect 180800 237134 181472 237218
rect 180800 236898 180858 237134
rect 181094 236898 181178 237134
rect 181414 236898 181472 237134
rect 180800 236866 181472 236898
rect 208000 237454 208672 237486
rect 208000 237218 208058 237454
rect 208294 237218 208378 237454
rect 208614 237218 208672 237454
rect 208000 237134 208672 237218
rect 208000 236898 208058 237134
rect 208294 236898 208378 237134
rect 208614 236898 208672 237134
rect 208000 236866 208672 236898
rect 235200 237454 235872 237486
rect 235200 237218 235258 237454
rect 235494 237218 235578 237454
rect 235814 237218 235872 237454
rect 235200 237134 235872 237218
rect 235200 236898 235258 237134
rect 235494 236898 235578 237134
rect 235814 236898 235872 237134
rect 235200 236866 235872 236898
rect 262400 237454 263072 237486
rect 262400 237218 262458 237454
rect 262694 237218 262778 237454
rect 263014 237218 263072 237454
rect 262400 237134 263072 237218
rect 262400 236898 262458 237134
rect 262694 236898 262778 237134
rect 263014 236898 263072 237134
rect 262400 236866 263072 236898
rect 289600 237454 290272 237486
rect 289600 237218 289658 237454
rect 289894 237218 289978 237454
rect 290214 237218 290272 237454
rect 289600 237134 290272 237218
rect 289600 236898 289658 237134
rect 289894 236898 289978 237134
rect 290214 236898 290272 237134
rect 289600 236866 290272 236898
rect 316800 237454 317472 237486
rect 316800 237218 316858 237454
rect 317094 237218 317178 237454
rect 317414 237218 317472 237454
rect 316800 237134 317472 237218
rect 316800 236898 316858 237134
rect 317094 236898 317178 237134
rect 317414 236898 317472 237134
rect 316800 236866 317472 236898
rect 344000 237454 344672 237486
rect 344000 237218 344058 237454
rect 344294 237218 344378 237454
rect 344614 237218 344672 237454
rect 344000 237134 344672 237218
rect 344000 236898 344058 237134
rect 344294 236898 344378 237134
rect 344614 236898 344672 237134
rect 344000 236866 344672 236898
rect 371200 237454 371872 237486
rect 371200 237218 371258 237454
rect 371494 237218 371578 237454
rect 371814 237218 371872 237454
rect 371200 237134 371872 237218
rect 371200 236898 371258 237134
rect 371494 236898 371578 237134
rect 371814 236898 371872 237134
rect 371200 236866 371872 236898
rect 398400 237454 399072 237486
rect 398400 237218 398458 237454
rect 398694 237218 398778 237454
rect 399014 237218 399072 237454
rect 398400 237134 399072 237218
rect 398400 236898 398458 237134
rect 398694 236898 398778 237134
rect 399014 236898 399072 237134
rect 398400 236866 399072 236898
rect 425600 237454 426272 237486
rect 425600 237218 425658 237454
rect 425894 237218 425978 237454
rect 426214 237218 426272 237454
rect 425600 237134 426272 237218
rect 425600 236898 425658 237134
rect 425894 236898 425978 237134
rect 426214 236898 426272 237134
rect 425600 236866 426272 236898
rect 452800 237454 453472 237486
rect 452800 237218 452858 237454
rect 453094 237218 453178 237454
rect 453414 237218 453472 237454
rect 452800 237134 453472 237218
rect 452800 236898 452858 237134
rect 453094 236898 453178 237134
rect 453414 236898 453472 237134
rect 452800 236866 453472 236898
rect 480000 237454 480672 237486
rect 480000 237218 480058 237454
rect 480294 237218 480378 237454
rect 480614 237218 480672 237454
rect 480000 237134 480672 237218
rect 480000 236898 480058 237134
rect 480294 236898 480378 237134
rect 480614 236898 480672 237134
rect 480000 236866 480672 236898
rect 507200 237454 507872 237486
rect 507200 237218 507258 237454
rect 507494 237218 507578 237454
rect 507814 237218 507872 237454
rect 507200 237134 507872 237218
rect 507200 236898 507258 237134
rect 507494 236898 507578 237134
rect 507814 236898 507872 237134
rect 507200 236866 507872 236898
rect 534400 237454 535072 237486
rect 534400 237218 534458 237454
rect 534694 237218 534778 237454
rect 535014 237218 535072 237454
rect 534400 237134 535072 237218
rect 534400 236898 534458 237134
rect 534694 236898 534778 237134
rect 535014 236898 535072 237134
rect 534400 236866 535072 236898
rect 561600 237454 562272 237486
rect 561600 237218 561658 237454
rect 561894 237218 561978 237454
rect 562214 237218 562272 237454
rect 561600 237134 562272 237218
rect 561600 236898 561658 237134
rect 561894 236898 561978 237134
rect 562214 236898 562272 237134
rect 561600 236866 562272 236898
rect 571500 237454 572120 237486
rect 571500 237218 571532 237454
rect 571768 237218 571852 237454
rect 572088 237218 572120 237454
rect 571500 237134 572120 237218
rect 571500 236898 571532 237134
rect 571768 236898 571852 237134
rect 572088 236898 572120 237134
rect 571500 236866 572120 236898
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect 9084 219454 9704 219486
rect 9084 219218 9116 219454
rect 9352 219218 9436 219454
rect 9672 219218 9704 219454
rect 9084 219134 9704 219218
rect 9084 218898 9116 219134
rect 9352 218898 9436 219134
rect 9672 218898 9704 219134
rect 9084 218866 9704 218898
rect 31200 219454 31872 219486
rect 31200 219218 31258 219454
rect 31494 219218 31578 219454
rect 31814 219218 31872 219454
rect 31200 219134 31872 219218
rect 31200 218898 31258 219134
rect 31494 218898 31578 219134
rect 31814 218898 31872 219134
rect 31200 218866 31872 218898
rect 35555 219454 35915 219486
rect 35555 219218 35617 219454
rect 35853 219218 35915 219454
rect 35555 219134 35915 219218
rect 35555 218898 35617 219134
rect 35853 218898 35915 219134
rect 35555 218866 35915 218898
rect 132591 219454 132951 219486
rect 132591 219218 132653 219454
rect 132889 219218 132951 219454
rect 132591 219134 132951 219218
rect 132591 218898 132653 219134
rect 132889 218898 132951 219134
rect 132591 218866 132951 218898
rect 139527 219454 139887 219486
rect 139527 219218 139589 219454
rect 139825 219218 139887 219454
rect 139527 219134 139887 219218
rect 139527 218898 139589 219134
rect 139825 218898 139887 219134
rect 139527 218866 139887 218898
rect 236563 219454 236923 219486
rect 236563 219218 236625 219454
rect 236861 219218 236923 219454
rect 236563 219134 236923 219218
rect 236563 218898 236625 219134
rect 236861 218898 236923 219134
rect 236563 218866 236923 218898
rect 248800 219454 249472 219486
rect 248800 219218 248858 219454
rect 249094 219218 249178 219454
rect 249414 219218 249472 219454
rect 248800 219134 249472 219218
rect 248800 218898 248858 219134
rect 249094 218898 249178 219134
rect 249414 218898 249472 219134
rect 248800 218866 249472 218898
rect 276000 219454 276672 219486
rect 276000 219218 276058 219454
rect 276294 219218 276378 219454
rect 276614 219218 276672 219454
rect 276000 219134 276672 219218
rect 276000 218898 276058 219134
rect 276294 218898 276378 219134
rect 276614 218898 276672 219134
rect 276000 218866 276672 218898
rect 303200 219454 303872 219486
rect 303200 219218 303258 219454
rect 303494 219218 303578 219454
rect 303814 219218 303872 219454
rect 303200 219134 303872 219218
rect 303200 218898 303258 219134
rect 303494 218898 303578 219134
rect 303814 218898 303872 219134
rect 303200 218866 303872 218898
rect 330400 219454 331072 219486
rect 330400 219218 330458 219454
rect 330694 219218 330778 219454
rect 331014 219218 331072 219454
rect 330400 219134 331072 219218
rect 330400 218898 330458 219134
rect 330694 218898 330778 219134
rect 331014 218898 331072 219134
rect 330400 218866 331072 218898
rect 342483 219454 342843 219486
rect 342483 219218 342545 219454
rect 342781 219218 342843 219454
rect 342483 219134 342843 219218
rect 342483 218898 342545 219134
rect 342781 218898 342843 219134
rect 342483 218866 342843 218898
rect 439519 219454 439879 219486
rect 439519 219218 439581 219454
rect 439817 219218 439879 219454
rect 439519 219134 439879 219218
rect 439519 218898 439581 219134
rect 439817 218898 439879 219134
rect 439519 218866 439879 218898
rect 446455 219454 446815 219486
rect 446455 219218 446517 219454
rect 446753 219218 446815 219454
rect 446455 219134 446815 219218
rect 446455 218898 446517 219134
rect 446753 218898 446815 219134
rect 446455 218866 446815 218898
rect 543491 219454 543851 219486
rect 543491 219218 543553 219454
rect 543789 219218 543851 219454
rect 543491 219134 543851 219218
rect 543491 218898 543553 219134
rect 543789 218898 543851 219134
rect 543491 218866 543851 218898
rect 548000 219454 548672 219486
rect 548000 219218 548058 219454
rect 548294 219218 548378 219454
rect 548614 219218 548672 219454
rect 548000 219134 548672 219218
rect 548000 218898 548058 219134
rect 548294 218898 548378 219134
rect 548614 218898 548672 219134
rect 548000 218866 548672 218898
rect 570260 219454 570880 219486
rect 570260 219218 570292 219454
rect 570528 219218 570612 219454
rect 570848 219218 570880 219454
rect 570260 219134 570880 219218
rect 570260 218898 570292 219134
rect 570528 218898 570612 219134
rect 570848 218898 570880 219134
rect 570260 218866 570880 218898
rect 7844 201454 8464 201486
rect 7844 201218 7876 201454
rect 8112 201218 8196 201454
rect 8432 201218 8464 201454
rect 7844 201134 8464 201218
rect 7844 200898 7876 201134
rect 8112 200898 8196 201134
rect 8432 200898 8464 201134
rect 7844 200866 8464 200898
rect 17600 201454 18272 201486
rect 17600 201218 17658 201454
rect 17894 201218 17978 201454
rect 18214 201218 18272 201454
rect 17600 201134 18272 201218
rect 17600 200898 17658 201134
rect 17894 200898 17978 201134
rect 18214 200898 18272 201134
rect 17600 200866 18272 200898
rect 34835 201454 35195 201486
rect 34835 201218 34897 201454
rect 35133 201218 35195 201454
rect 34835 201134 35195 201218
rect 34835 200898 34897 201134
rect 35133 200898 35195 201134
rect 34835 200866 35195 200898
rect 133311 201454 133671 201486
rect 133311 201218 133373 201454
rect 133609 201218 133671 201454
rect 133311 201134 133671 201218
rect 133311 200898 133373 201134
rect 133609 200898 133671 201134
rect 133311 200866 133671 200898
rect 138807 201454 139167 201486
rect 138807 201218 138869 201454
rect 139105 201218 139167 201454
rect 138807 201134 139167 201218
rect 138807 200898 138869 201134
rect 139105 200898 139167 201134
rect 138807 200866 139167 200898
rect 237283 201454 237643 201486
rect 237283 201218 237345 201454
rect 237581 201218 237643 201454
rect 237283 201134 237643 201218
rect 237283 200898 237345 201134
rect 237581 200898 237643 201134
rect 237283 200866 237643 200898
rect 262400 201454 263072 201486
rect 262400 201218 262458 201454
rect 262694 201218 262778 201454
rect 263014 201218 263072 201454
rect 262400 201134 263072 201218
rect 262400 200898 262458 201134
rect 262694 200898 262778 201134
rect 263014 200898 263072 201134
rect 262400 200866 263072 200898
rect 289600 201454 290272 201486
rect 289600 201218 289658 201454
rect 289894 201218 289978 201454
rect 290214 201218 290272 201454
rect 289600 201134 290272 201218
rect 289600 200898 289658 201134
rect 289894 200898 289978 201134
rect 290214 200898 290272 201134
rect 289600 200866 290272 200898
rect 316800 201454 317472 201486
rect 316800 201218 316858 201454
rect 317094 201218 317178 201454
rect 317414 201218 317472 201454
rect 316800 201134 317472 201218
rect 316800 200898 316858 201134
rect 317094 200898 317178 201134
rect 317414 200898 317472 201134
rect 316800 200866 317472 200898
rect 341763 201454 342123 201486
rect 341763 201218 341825 201454
rect 342061 201218 342123 201454
rect 341763 201134 342123 201218
rect 341763 200898 341825 201134
rect 342061 200898 342123 201134
rect 341763 200866 342123 200898
rect 440239 201454 440599 201486
rect 440239 201218 440301 201454
rect 440537 201218 440599 201454
rect 440239 201134 440599 201218
rect 440239 200898 440301 201134
rect 440537 200898 440599 201134
rect 440239 200866 440599 200898
rect 445735 201454 446095 201486
rect 445735 201218 445797 201454
rect 446033 201218 446095 201454
rect 445735 201134 446095 201218
rect 445735 200898 445797 201134
rect 446033 200898 446095 201134
rect 445735 200866 446095 200898
rect 544211 201454 544571 201486
rect 544211 201218 544273 201454
rect 544509 201218 544571 201454
rect 544211 201134 544571 201218
rect 544211 200898 544273 201134
rect 544509 200898 544571 201134
rect 544211 200866 544571 200898
rect 561600 201454 562272 201486
rect 561600 201218 561658 201454
rect 561894 201218 561978 201454
rect 562214 201218 562272 201454
rect 561600 201134 562272 201218
rect 561600 200898 561658 201134
rect 561894 200898 561978 201134
rect 562214 200898 562272 201134
rect 561600 200866 562272 200898
rect 571500 201454 572120 201486
rect 571500 201218 571532 201454
rect 571768 201218 571852 201454
rect 572088 201218 572120 201454
rect 571500 201134 572120 201218
rect 571500 200898 571532 201134
rect 571768 200898 571852 201134
rect 572088 200898 572120 201134
rect 571500 200866 572120 200898
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect 9084 183454 9704 183486
rect 9084 183218 9116 183454
rect 9352 183218 9436 183454
rect 9672 183218 9704 183454
rect 9084 183134 9704 183218
rect 9084 182898 9116 183134
rect 9352 182898 9436 183134
rect 9672 182898 9704 183134
rect 9084 182866 9704 182898
rect 31200 183454 31872 183486
rect 31200 183218 31258 183454
rect 31494 183218 31578 183454
rect 31814 183218 31872 183454
rect 31200 183134 31872 183218
rect 31200 182898 31258 183134
rect 31494 182898 31578 183134
rect 31814 182898 31872 183134
rect 31200 182866 31872 182898
rect 35555 183454 35915 183486
rect 35555 183218 35617 183454
rect 35853 183218 35915 183454
rect 35555 183134 35915 183218
rect 35555 182898 35617 183134
rect 35853 182898 35915 183134
rect 35555 182866 35915 182898
rect 132591 183454 132951 183486
rect 132591 183218 132653 183454
rect 132889 183218 132951 183454
rect 132591 183134 132951 183218
rect 132591 182898 132653 183134
rect 132889 182898 132951 183134
rect 132591 182866 132951 182898
rect 139527 183454 139887 183486
rect 139527 183218 139589 183454
rect 139825 183218 139887 183454
rect 139527 183134 139887 183218
rect 139527 182898 139589 183134
rect 139825 182898 139887 183134
rect 139527 182866 139887 182898
rect 236563 183454 236923 183486
rect 236563 183218 236625 183454
rect 236861 183218 236923 183454
rect 236563 183134 236923 183218
rect 236563 182898 236625 183134
rect 236861 182898 236923 183134
rect 236563 182866 236923 182898
rect 248800 183454 249472 183486
rect 248800 183218 248858 183454
rect 249094 183218 249178 183454
rect 249414 183218 249472 183454
rect 248800 183134 249472 183218
rect 248800 182898 248858 183134
rect 249094 182898 249178 183134
rect 249414 182898 249472 183134
rect 248800 182866 249472 182898
rect 276000 183454 276672 183486
rect 276000 183218 276058 183454
rect 276294 183218 276378 183454
rect 276614 183218 276672 183454
rect 276000 183134 276672 183218
rect 276000 182898 276058 183134
rect 276294 182898 276378 183134
rect 276614 182898 276672 183134
rect 276000 182866 276672 182898
rect 303200 183454 303872 183486
rect 303200 183218 303258 183454
rect 303494 183218 303578 183454
rect 303814 183218 303872 183454
rect 303200 183134 303872 183218
rect 303200 182898 303258 183134
rect 303494 182898 303578 183134
rect 303814 182898 303872 183134
rect 303200 182866 303872 182898
rect 330400 183454 331072 183486
rect 330400 183218 330458 183454
rect 330694 183218 330778 183454
rect 331014 183218 331072 183454
rect 330400 183134 331072 183218
rect 330400 182898 330458 183134
rect 330694 182898 330778 183134
rect 331014 182898 331072 183134
rect 330400 182866 331072 182898
rect 342483 183454 342843 183486
rect 342483 183218 342545 183454
rect 342781 183218 342843 183454
rect 342483 183134 342843 183218
rect 342483 182898 342545 183134
rect 342781 182898 342843 183134
rect 342483 182866 342843 182898
rect 439519 183454 439879 183486
rect 439519 183218 439581 183454
rect 439817 183218 439879 183454
rect 439519 183134 439879 183218
rect 439519 182898 439581 183134
rect 439817 182898 439879 183134
rect 439519 182866 439879 182898
rect 446455 183454 446815 183486
rect 446455 183218 446517 183454
rect 446753 183218 446815 183454
rect 446455 183134 446815 183218
rect 446455 182898 446517 183134
rect 446753 182898 446815 183134
rect 446455 182866 446815 182898
rect 543491 183454 543851 183486
rect 543491 183218 543553 183454
rect 543789 183218 543851 183454
rect 543491 183134 543851 183218
rect 543491 182898 543553 183134
rect 543789 182898 543851 183134
rect 543491 182866 543851 182898
rect 548000 183454 548672 183486
rect 548000 183218 548058 183454
rect 548294 183218 548378 183454
rect 548614 183218 548672 183454
rect 548000 183134 548672 183218
rect 548000 182898 548058 183134
rect 548294 182898 548378 183134
rect 548614 182898 548672 183134
rect 548000 182866 548672 182898
rect 570260 183454 570880 183486
rect 570260 183218 570292 183454
rect 570528 183218 570612 183454
rect 570848 183218 570880 183454
rect 570260 183134 570880 183218
rect 570260 182898 570292 183134
rect 570528 182898 570612 183134
rect 570848 182898 570880 183134
rect 570260 182866 570880 182898
rect 7844 165454 8464 165486
rect 7844 165218 7876 165454
rect 8112 165218 8196 165454
rect 8432 165218 8464 165454
rect 7844 165134 8464 165218
rect 7844 164898 7876 165134
rect 8112 164898 8196 165134
rect 8432 164898 8464 165134
rect 7844 164866 8464 164898
rect 17600 165454 18272 165486
rect 17600 165218 17658 165454
rect 17894 165218 17978 165454
rect 18214 165218 18272 165454
rect 17600 165134 18272 165218
rect 17600 164898 17658 165134
rect 17894 164898 17978 165134
rect 18214 164898 18272 165134
rect 17600 164866 18272 164898
rect 34835 165454 35195 165486
rect 34835 165218 34897 165454
rect 35133 165218 35195 165454
rect 34835 165134 35195 165218
rect 34835 164898 34897 165134
rect 35133 164898 35195 165134
rect 34835 164866 35195 164898
rect 133311 165454 133671 165486
rect 133311 165218 133373 165454
rect 133609 165218 133671 165454
rect 133311 165134 133671 165218
rect 133311 164898 133373 165134
rect 133609 164898 133671 165134
rect 133311 164866 133671 164898
rect 138807 165454 139167 165486
rect 138807 165218 138869 165454
rect 139105 165218 139167 165454
rect 138807 165134 139167 165218
rect 138807 164898 138869 165134
rect 139105 164898 139167 165134
rect 138807 164866 139167 164898
rect 237283 165454 237643 165486
rect 237283 165218 237345 165454
rect 237581 165218 237643 165454
rect 237283 165134 237643 165218
rect 237283 164898 237345 165134
rect 237581 164898 237643 165134
rect 237283 164866 237643 164898
rect 262400 165454 263072 165486
rect 262400 165218 262458 165454
rect 262694 165218 262778 165454
rect 263014 165218 263072 165454
rect 262400 165134 263072 165218
rect 262400 164898 262458 165134
rect 262694 164898 262778 165134
rect 263014 164898 263072 165134
rect 262400 164866 263072 164898
rect 289600 165454 290272 165486
rect 289600 165218 289658 165454
rect 289894 165218 289978 165454
rect 290214 165218 290272 165454
rect 289600 165134 290272 165218
rect 289600 164898 289658 165134
rect 289894 164898 289978 165134
rect 290214 164898 290272 165134
rect 289600 164866 290272 164898
rect 316800 165454 317472 165486
rect 316800 165218 316858 165454
rect 317094 165218 317178 165454
rect 317414 165218 317472 165454
rect 316800 165134 317472 165218
rect 316800 164898 316858 165134
rect 317094 164898 317178 165134
rect 317414 164898 317472 165134
rect 316800 164866 317472 164898
rect 341763 165454 342123 165486
rect 341763 165218 341825 165454
rect 342061 165218 342123 165454
rect 341763 165134 342123 165218
rect 341763 164898 341825 165134
rect 342061 164898 342123 165134
rect 341763 164866 342123 164898
rect 440239 165454 440599 165486
rect 440239 165218 440301 165454
rect 440537 165218 440599 165454
rect 440239 165134 440599 165218
rect 440239 164898 440301 165134
rect 440537 164898 440599 165134
rect 440239 164866 440599 164898
rect 445735 165454 446095 165486
rect 445735 165218 445797 165454
rect 446033 165218 446095 165454
rect 445735 165134 446095 165218
rect 445735 164898 445797 165134
rect 446033 164898 446095 165134
rect 445735 164866 446095 164898
rect 544211 165454 544571 165486
rect 544211 165218 544273 165454
rect 544509 165218 544571 165454
rect 544211 165134 544571 165218
rect 544211 164898 544273 165134
rect 544509 164898 544571 165134
rect 544211 164866 544571 164898
rect 561600 165454 562272 165486
rect 561600 165218 561658 165454
rect 561894 165218 561978 165454
rect 562214 165218 562272 165454
rect 561600 165134 562272 165218
rect 561600 164898 561658 165134
rect 561894 164898 561978 165134
rect 562214 164898 562272 165134
rect 561600 164866 562272 164898
rect 571500 165454 572120 165486
rect 571500 165218 571532 165454
rect 571768 165218 571852 165454
rect 572088 165218 572120 165454
rect 571500 165134 572120 165218
rect 571500 164898 571532 165134
rect 571768 164898 571852 165134
rect 572088 164898 572120 165134
rect 571500 164866 572120 164898
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect 9084 147454 9704 147486
rect 9084 147218 9116 147454
rect 9352 147218 9436 147454
rect 9672 147218 9704 147454
rect 9084 147134 9704 147218
rect 9084 146898 9116 147134
rect 9352 146898 9436 147134
rect 9672 146898 9704 147134
rect 9084 146866 9704 146898
rect 31200 147454 31872 147486
rect 31200 147218 31258 147454
rect 31494 147218 31578 147454
rect 31814 147218 31872 147454
rect 31200 147134 31872 147218
rect 31200 146898 31258 147134
rect 31494 146898 31578 147134
rect 31814 146898 31872 147134
rect 31200 146866 31872 146898
rect 58400 147454 59072 147486
rect 58400 147218 58458 147454
rect 58694 147218 58778 147454
rect 59014 147218 59072 147454
rect 58400 147134 59072 147218
rect 58400 146898 58458 147134
rect 58694 146898 58778 147134
rect 59014 146898 59072 147134
rect 58400 146866 59072 146898
rect 85600 147454 86272 147486
rect 85600 147218 85658 147454
rect 85894 147218 85978 147454
rect 86214 147218 86272 147454
rect 85600 147134 86272 147218
rect 85600 146898 85658 147134
rect 85894 146898 85978 147134
rect 86214 146898 86272 147134
rect 85600 146866 86272 146898
rect 112800 147454 113472 147486
rect 112800 147218 112858 147454
rect 113094 147218 113178 147454
rect 113414 147218 113472 147454
rect 112800 147134 113472 147218
rect 112800 146898 112858 147134
rect 113094 146898 113178 147134
rect 113414 146898 113472 147134
rect 112800 146866 113472 146898
rect 140000 147454 140672 147486
rect 140000 147218 140058 147454
rect 140294 147218 140378 147454
rect 140614 147218 140672 147454
rect 140000 147134 140672 147218
rect 140000 146898 140058 147134
rect 140294 146898 140378 147134
rect 140614 146898 140672 147134
rect 140000 146866 140672 146898
rect 167200 147454 167872 147486
rect 167200 147218 167258 147454
rect 167494 147218 167578 147454
rect 167814 147218 167872 147454
rect 167200 147134 167872 147218
rect 167200 146898 167258 147134
rect 167494 146898 167578 147134
rect 167814 146898 167872 147134
rect 167200 146866 167872 146898
rect 194400 147454 195072 147486
rect 194400 147218 194458 147454
rect 194694 147218 194778 147454
rect 195014 147218 195072 147454
rect 194400 147134 195072 147218
rect 194400 146898 194458 147134
rect 194694 146898 194778 147134
rect 195014 146898 195072 147134
rect 194400 146866 195072 146898
rect 221600 147454 222272 147486
rect 221600 147218 221658 147454
rect 221894 147218 221978 147454
rect 222214 147218 222272 147454
rect 221600 147134 222272 147218
rect 221600 146898 221658 147134
rect 221894 146898 221978 147134
rect 222214 146898 222272 147134
rect 221600 146866 222272 146898
rect 248800 147454 249472 147486
rect 248800 147218 248858 147454
rect 249094 147218 249178 147454
rect 249414 147218 249472 147454
rect 248800 147134 249472 147218
rect 248800 146898 248858 147134
rect 249094 146898 249178 147134
rect 249414 146898 249472 147134
rect 248800 146866 249472 146898
rect 276000 147454 276672 147486
rect 276000 147218 276058 147454
rect 276294 147218 276378 147454
rect 276614 147218 276672 147454
rect 276000 147134 276672 147218
rect 276000 146898 276058 147134
rect 276294 146898 276378 147134
rect 276614 146898 276672 147134
rect 276000 146866 276672 146898
rect 303200 147454 303872 147486
rect 303200 147218 303258 147454
rect 303494 147218 303578 147454
rect 303814 147218 303872 147454
rect 303200 147134 303872 147218
rect 303200 146898 303258 147134
rect 303494 146898 303578 147134
rect 303814 146898 303872 147134
rect 303200 146866 303872 146898
rect 330400 147454 331072 147486
rect 330400 147218 330458 147454
rect 330694 147218 330778 147454
rect 331014 147218 331072 147454
rect 330400 147134 331072 147218
rect 330400 146898 330458 147134
rect 330694 146898 330778 147134
rect 331014 146898 331072 147134
rect 330400 146866 331072 146898
rect 357600 147454 358272 147486
rect 357600 147218 357658 147454
rect 357894 147218 357978 147454
rect 358214 147218 358272 147454
rect 357600 147134 358272 147218
rect 357600 146898 357658 147134
rect 357894 146898 357978 147134
rect 358214 146898 358272 147134
rect 357600 146866 358272 146898
rect 384800 147454 385472 147486
rect 384800 147218 384858 147454
rect 385094 147218 385178 147454
rect 385414 147218 385472 147454
rect 384800 147134 385472 147218
rect 384800 146898 384858 147134
rect 385094 146898 385178 147134
rect 385414 146898 385472 147134
rect 384800 146866 385472 146898
rect 412000 147454 412672 147486
rect 412000 147218 412058 147454
rect 412294 147218 412378 147454
rect 412614 147218 412672 147454
rect 412000 147134 412672 147218
rect 412000 146898 412058 147134
rect 412294 146898 412378 147134
rect 412614 146898 412672 147134
rect 412000 146866 412672 146898
rect 439200 147454 439872 147486
rect 439200 147218 439258 147454
rect 439494 147218 439578 147454
rect 439814 147218 439872 147454
rect 439200 147134 439872 147218
rect 439200 146898 439258 147134
rect 439494 146898 439578 147134
rect 439814 146898 439872 147134
rect 439200 146866 439872 146898
rect 466400 147454 467072 147486
rect 466400 147218 466458 147454
rect 466694 147218 466778 147454
rect 467014 147218 467072 147454
rect 466400 147134 467072 147218
rect 466400 146898 466458 147134
rect 466694 146898 466778 147134
rect 467014 146898 467072 147134
rect 466400 146866 467072 146898
rect 493600 147454 494272 147486
rect 493600 147218 493658 147454
rect 493894 147218 493978 147454
rect 494214 147218 494272 147454
rect 493600 147134 494272 147218
rect 493600 146898 493658 147134
rect 493894 146898 493978 147134
rect 494214 146898 494272 147134
rect 493600 146866 494272 146898
rect 520800 147454 521472 147486
rect 520800 147218 520858 147454
rect 521094 147218 521178 147454
rect 521414 147218 521472 147454
rect 520800 147134 521472 147218
rect 520800 146898 520858 147134
rect 521094 146898 521178 147134
rect 521414 146898 521472 147134
rect 520800 146866 521472 146898
rect 548000 147454 548672 147486
rect 548000 147218 548058 147454
rect 548294 147218 548378 147454
rect 548614 147218 548672 147454
rect 548000 147134 548672 147218
rect 548000 146898 548058 147134
rect 548294 146898 548378 147134
rect 548614 146898 548672 147134
rect 548000 146866 548672 146898
rect 570260 147454 570880 147486
rect 570260 147218 570292 147454
rect 570528 147218 570612 147454
rect 570848 147218 570880 147454
rect 570260 147134 570880 147218
rect 570260 146898 570292 147134
rect 570528 146898 570612 147134
rect 570848 146898 570880 147134
rect 570260 146866 570880 146898
rect 7844 129454 8464 129486
rect 7844 129218 7876 129454
rect 8112 129218 8196 129454
rect 8432 129218 8464 129454
rect 7844 129134 8464 129218
rect 7844 128898 7876 129134
rect 8112 128898 8196 129134
rect 8432 128898 8464 129134
rect 7844 128866 8464 128898
rect 17600 129454 18272 129486
rect 17600 129218 17658 129454
rect 17894 129218 17978 129454
rect 18214 129218 18272 129454
rect 17600 129134 18272 129218
rect 17600 128898 17658 129134
rect 17894 128898 17978 129134
rect 18214 128898 18272 129134
rect 17600 128866 18272 128898
rect 34835 129454 35195 129486
rect 34835 129218 34897 129454
rect 35133 129218 35195 129454
rect 34835 129134 35195 129218
rect 34835 128898 34897 129134
rect 35133 128898 35195 129134
rect 34835 128866 35195 128898
rect 133311 129454 133671 129486
rect 133311 129218 133373 129454
rect 133609 129218 133671 129454
rect 133311 129134 133671 129218
rect 133311 128898 133373 129134
rect 133609 128898 133671 129134
rect 133311 128866 133671 128898
rect 138807 129454 139167 129486
rect 138807 129218 138869 129454
rect 139105 129218 139167 129454
rect 138807 129134 139167 129218
rect 138807 128898 138869 129134
rect 139105 128898 139167 129134
rect 138807 128866 139167 128898
rect 237283 129454 237643 129486
rect 237283 129218 237345 129454
rect 237581 129218 237643 129454
rect 237283 129134 237643 129218
rect 237283 128898 237345 129134
rect 237581 128898 237643 129134
rect 237283 128866 237643 128898
rect 262400 129454 263072 129486
rect 262400 129218 262458 129454
rect 262694 129218 262778 129454
rect 263014 129218 263072 129454
rect 262400 129134 263072 129218
rect 262400 128898 262458 129134
rect 262694 128898 262778 129134
rect 263014 128898 263072 129134
rect 262400 128866 263072 128898
rect 289600 129454 290272 129486
rect 289600 129218 289658 129454
rect 289894 129218 289978 129454
rect 290214 129218 290272 129454
rect 289600 129134 290272 129218
rect 289600 128898 289658 129134
rect 289894 128898 289978 129134
rect 290214 128898 290272 129134
rect 289600 128866 290272 128898
rect 316800 129454 317472 129486
rect 316800 129218 316858 129454
rect 317094 129218 317178 129454
rect 317414 129218 317472 129454
rect 316800 129134 317472 129218
rect 316800 128898 316858 129134
rect 317094 128898 317178 129134
rect 317414 128898 317472 129134
rect 316800 128866 317472 128898
rect 341763 129454 342123 129486
rect 341763 129218 341825 129454
rect 342061 129218 342123 129454
rect 341763 129134 342123 129218
rect 341763 128898 341825 129134
rect 342061 128898 342123 129134
rect 341763 128866 342123 128898
rect 440239 129454 440599 129486
rect 440239 129218 440301 129454
rect 440537 129218 440599 129454
rect 440239 129134 440599 129218
rect 440239 128898 440301 129134
rect 440537 128898 440599 129134
rect 440239 128866 440599 128898
rect 445735 129454 446095 129486
rect 445735 129218 445797 129454
rect 446033 129218 446095 129454
rect 445735 129134 446095 129218
rect 445735 128898 445797 129134
rect 446033 128898 446095 129134
rect 445735 128866 446095 128898
rect 544211 129454 544571 129486
rect 544211 129218 544273 129454
rect 544509 129218 544571 129454
rect 544211 129134 544571 129218
rect 544211 128898 544273 129134
rect 544509 128898 544571 129134
rect 544211 128866 544571 128898
rect 561600 129454 562272 129486
rect 561600 129218 561658 129454
rect 561894 129218 561978 129454
rect 562214 129218 562272 129454
rect 561600 129134 562272 129218
rect 561600 128898 561658 129134
rect 561894 128898 561978 129134
rect 562214 128898 562272 129134
rect 561600 128866 562272 128898
rect 571500 129454 572120 129486
rect 571500 129218 571532 129454
rect 571768 129218 571852 129454
rect 572088 129218 572120 129454
rect 571500 129134 572120 129218
rect 571500 128898 571532 129134
rect 571768 128898 571852 129134
rect 572088 128898 572120 129134
rect 571500 128866 572120 128898
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect 9084 111454 9704 111486
rect 9084 111218 9116 111454
rect 9352 111218 9436 111454
rect 9672 111218 9704 111454
rect 9084 111134 9704 111218
rect 9084 110898 9116 111134
rect 9352 110898 9436 111134
rect 9672 110898 9704 111134
rect 9084 110866 9704 110898
rect 31200 111454 31872 111486
rect 31200 111218 31258 111454
rect 31494 111218 31578 111454
rect 31814 111218 31872 111454
rect 31200 111134 31872 111218
rect 31200 110898 31258 111134
rect 31494 110898 31578 111134
rect 31814 110898 31872 111134
rect 31200 110866 31872 110898
rect 35555 111454 35915 111486
rect 35555 111218 35617 111454
rect 35853 111218 35915 111454
rect 35555 111134 35915 111218
rect 35555 110898 35617 111134
rect 35853 110898 35915 111134
rect 35555 110866 35915 110898
rect 132591 111454 132951 111486
rect 132591 111218 132653 111454
rect 132889 111218 132951 111454
rect 132591 111134 132951 111218
rect 132591 110898 132653 111134
rect 132889 110898 132951 111134
rect 132591 110866 132951 110898
rect 139527 111454 139887 111486
rect 139527 111218 139589 111454
rect 139825 111218 139887 111454
rect 139527 111134 139887 111218
rect 139527 110898 139589 111134
rect 139825 110898 139887 111134
rect 139527 110866 139887 110898
rect 236563 111454 236923 111486
rect 236563 111218 236625 111454
rect 236861 111218 236923 111454
rect 236563 111134 236923 111218
rect 236563 110898 236625 111134
rect 236861 110898 236923 111134
rect 236563 110866 236923 110898
rect 248800 111454 249472 111486
rect 248800 111218 248858 111454
rect 249094 111218 249178 111454
rect 249414 111218 249472 111454
rect 248800 111134 249472 111218
rect 248800 110898 248858 111134
rect 249094 110898 249178 111134
rect 249414 110898 249472 111134
rect 248800 110866 249472 110898
rect 276000 111454 276672 111486
rect 276000 111218 276058 111454
rect 276294 111218 276378 111454
rect 276614 111218 276672 111454
rect 276000 111134 276672 111218
rect 276000 110898 276058 111134
rect 276294 110898 276378 111134
rect 276614 110898 276672 111134
rect 276000 110866 276672 110898
rect 303200 111454 303872 111486
rect 303200 111218 303258 111454
rect 303494 111218 303578 111454
rect 303814 111218 303872 111454
rect 303200 111134 303872 111218
rect 303200 110898 303258 111134
rect 303494 110898 303578 111134
rect 303814 110898 303872 111134
rect 303200 110866 303872 110898
rect 330400 111454 331072 111486
rect 330400 111218 330458 111454
rect 330694 111218 330778 111454
rect 331014 111218 331072 111454
rect 330400 111134 331072 111218
rect 330400 110898 330458 111134
rect 330694 110898 330778 111134
rect 331014 110898 331072 111134
rect 330400 110866 331072 110898
rect 342483 111454 342843 111486
rect 342483 111218 342545 111454
rect 342781 111218 342843 111454
rect 342483 111134 342843 111218
rect 342483 110898 342545 111134
rect 342781 110898 342843 111134
rect 342483 110866 342843 110898
rect 439519 111454 439879 111486
rect 439519 111218 439581 111454
rect 439817 111218 439879 111454
rect 439519 111134 439879 111218
rect 439519 110898 439581 111134
rect 439817 110898 439879 111134
rect 439519 110866 439879 110898
rect 446455 111454 446815 111486
rect 446455 111218 446517 111454
rect 446753 111218 446815 111454
rect 446455 111134 446815 111218
rect 446455 110898 446517 111134
rect 446753 110898 446815 111134
rect 446455 110866 446815 110898
rect 543491 111454 543851 111486
rect 543491 111218 543553 111454
rect 543789 111218 543851 111454
rect 543491 111134 543851 111218
rect 543491 110898 543553 111134
rect 543789 110898 543851 111134
rect 543491 110866 543851 110898
rect 548000 111454 548672 111486
rect 548000 111218 548058 111454
rect 548294 111218 548378 111454
rect 548614 111218 548672 111454
rect 548000 111134 548672 111218
rect 548000 110898 548058 111134
rect 548294 110898 548378 111134
rect 548614 110898 548672 111134
rect 548000 110866 548672 110898
rect 570260 111454 570880 111486
rect 570260 111218 570292 111454
rect 570528 111218 570612 111454
rect 570848 111218 570880 111454
rect 570260 111134 570880 111218
rect 570260 110898 570292 111134
rect 570528 110898 570612 111134
rect 570848 110898 570880 111134
rect 570260 110866 570880 110898
rect 7844 93454 8464 93486
rect 7844 93218 7876 93454
rect 8112 93218 8196 93454
rect 8432 93218 8464 93454
rect 7844 93134 8464 93218
rect 7844 92898 7876 93134
rect 8112 92898 8196 93134
rect 8432 92898 8464 93134
rect 7844 92866 8464 92898
rect 17600 93454 18272 93486
rect 17600 93218 17658 93454
rect 17894 93218 17978 93454
rect 18214 93218 18272 93454
rect 17600 93134 18272 93218
rect 17600 92898 17658 93134
rect 17894 92898 17978 93134
rect 18214 92898 18272 93134
rect 17600 92866 18272 92898
rect 34835 93454 35195 93486
rect 34835 93218 34897 93454
rect 35133 93218 35195 93454
rect 34835 93134 35195 93218
rect 34835 92898 34897 93134
rect 35133 92898 35195 93134
rect 34835 92866 35195 92898
rect 133311 93454 133671 93486
rect 133311 93218 133373 93454
rect 133609 93218 133671 93454
rect 133311 93134 133671 93218
rect 133311 92898 133373 93134
rect 133609 92898 133671 93134
rect 133311 92866 133671 92898
rect 138807 93454 139167 93486
rect 138807 93218 138869 93454
rect 139105 93218 139167 93454
rect 138807 93134 139167 93218
rect 138807 92898 138869 93134
rect 139105 92898 139167 93134
rect 138807 92866 139167 92898
rect 237283 93454 237643 93486
rect 237283 93218 237345 93454
rect 237581 93218 237643 93454
rect 237283 93134 237643 93218
rect 237283 92898 237345 93134
rect 237581 92898 237643 93134
rect 237283 92866 237643 92898
rect 262400 93454 263072 93486
rect 262400 93218 262458 93454
rect 262694 93218 262778 93454
rect 263014 93218 263072 93454
rect 262400 93134 263072 93218
rect 262400 92898 262458 93134
rect 262694 92898 262778 93134
rect 263014 92898 263072 93134
rect 262400 92866 263072 92898
rect 289600 93454 290272 93486
rect 289600 93218 289658 93454
rect 289894 93218 289978 93454
rect 290214 93218 290272 93454
rect 289600 93134 290272 93218
rect 289600 92898 289658 93134
rect 289894 92898 289978 93134
rect 290214 92898 290272 93134
rect 289600 92866 290272 92898
rect 316800 93454 317472 93486
rect 316800 93218 316858 93454
rect 317094 93218 317178 93454
rect 317414 93218 317472 93454
rect 316800 93134 317472 93218
rect 316800 92898 316858 93134
rect 317094 92898 317178 93134
rect 317414 92898 317472 93134
rect 316800 92866 317472 92898
rect 341763 93454 342123 93486
rect 341763 93218 341825 93454
rect 342061 93218 342123 93454
rect 341763 93134 342123 93218
rect 341763 92898 341825 93134
rect 342061 92898 342123 93134
rect 341763 92866 342123 92898
rect 440239 93454 440599 93486
rect 440239 93218 440301 93454
rect 440537 93218 440599 93454
rect 440239 93134 440599 93218
rect 440239 92898 440301 93134
rect 440537 92898 440599 93134
rect 440239 92866 440599 92898
rect 445735 93454 446095 93486
rect 445735 93218 445797 93454
rect 446033 93218 446095 93454
rect 445735 93134 446095 93218
rect 445735 92898 445797 93134
rect 446033 92898 446095 93134
rect 445735 92866 446095 92898
rect 544211 93454 544571 93486
rect 544211 93218 544273 93454
rect 544509 93218 544571 93454
rect 544211 93134 544571 93218
rect 544211 92898 544273 93134
rect 544509 92898 544571 93134
rect 544211 92866 544571 92898
rect 561600 93454 562272 93486
rect 561600 93218 561658 93454
rect 561894 93218 561978 93454
rect 562214 93218 562272 93454
rect 561600 93134 562272 93218
rect 561600 92898 561658 93134
rect 561894 92898 561978 93134
rect 562214 92898 562272 93134
rect 561600 92866 562272 92898
rect 571500 93454 572120 93486
rect 571500 93218 571532 93454
rect 571768 93218 571852 93454
rect 572088 93218 572120 93454
rect 571500 93134 572120 93218
rect 571500 92898 571532 93134
rect 571768 92898 571852 93134
rect 572088 92898 572120 93134
rect 571500 92866 572120 92898
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect 9084 75454 9704 75486
rect 9084 75218 9116 75454
rect 9352 75218 9436 75454
rect 9672 75218 9704 75454
rect 9084 75134 9704 75218
rect 9084 74898 9116 75134
rect 9352 74898 9436 75134
rect 9672 74898 9704 75134
rect 9084 74866 9704 74898
rect 31200 75454 31872 75486
rect 31200 75218 31258 75454
rect 31494 75218 31578 75454
rect 31814 75218 31872 75454
rect 31200 75134 31872 75218
rect 31200 74898 31258 75134
rect 31494 74898 31578 75134
rect 31814 74898 31872 75134
rect 31200 74866 31872 74898
rect 35555 75454 35915 75486
rect 35555 75218 35617 75454
rect 35853 75218 35915 75454
rect 35555 75134 35915 75218
rect 35555 74898 35617 75134
rect 35853 74898 35915 75134
rect 35555 74866 35915 74898
rect 132591 75454 132951 75486
rect 132591 75218 132653 75454
rect 132889 75218 132951 75454
rect 132591 75134 132951 75218
rect 132591 74898 132653 75134
rect 132889 74898 132951 75134
rect 132591 74866 132951 74898
rect 139527 75454 139887 75486
rect 139527 75218 139589 75454
rect 139825 75218 139887 75454
rect 139527 75134 139887 75218
rect 139527 74898 139589 75134
rect 139825 74898 139887 75134
rect 139527 74866 139887 74898
rect 236563 75454 236923 75486
rect 236563 75218 236625 75454
rect 236861 75218 236923 75454
rect 236563 75134 236923 75218
rect 236563 74898 236625 75134
rect 236861 74898 236923 75134
rect 236563 74866 236923 74898
rect 248800 75454 249472 75486
rect 248800 75218 248858 75454
rect 249094 75218 249178 75454
rect 249414 75218 249472 75454
rect 248800 75134 249472 75218
rect 248800 74898 248858 75134
rect 249094 74898 249178 75134
rect 249414 74898 249472 75134
rect 248800 74866 249472 74898
rect 276000 75454 276672 75486
rect 276000 75218 276058 75454
rect 276294 75218 276378 75454
rect 276614 75218 276672 75454
rect 276000 75134 276672 75218
rect 276000 74898 276058 75134
rect 276294 74898 276378 75134
rect 276614 74898 276672 75134
rect 276000 74866 276672 74898
rect 303200 75454 303872 75486
rect 303200 75218 303258 75454
rect 303494 75218 303578 75454
rect 303814 75218 303872 75454
rect 303200 75134 303872 75218
rect 303200 74898 303258 75134
rect 303494 74898 303578 75134
rect 303814 74898 303872 75134
rect 303200 74866 303872 74898
rect 330400 75454 331072 75486
rect 330400 75218 330458 75454
rect 330694 75218 330778 75454
rect 331014 75218 331072 75454
rect 330400 75134 331072 75218
rect 330400 74898 330458 75134
rect 330694 74898 330778 75134
rect 331014 74898 331072 75134
rect 330400 74866 331072 74898
rect 342483 75454 342843 75486
rect 342483 75218 342545 75454
rect 342781 75218 342843 75454
rect 342483 75134 342843 75218
rect 342483 74898 342545 75134
rect 342781 74898 342843 75134
rect 342483 74866 342843 74898
rect 439519 75454 439879 75486
rect 439519 75218 439581 75454
rect 439817 75218 439879 75454
rect 439519 75134 439879 75218
rect 439519 74898 439581 75134
rect 439817 74898 439879 75134
rect 439519 74866 439879 74898
rect 446455 75454 446815 75486
rect 446455 75218 446517 75454
rect 446753 75218 446815 75454
rect 446455 75134 446815 75218
rect 446455 74898 446517 75134
rect 446753 74898 446815 75134
rect 446455 74866 446815 74898
rect 543491 75454 543851 75486
rect 543491 75218 543553 75454
rect 543789 75218 543851 75454
rect 543491 75134 543851 75218
rect 543491 74898 543553 75134
rect 543789 74898 543851 75134
rect 543491 74866 543851 74898
rect 548000 75454 548672 75486
rect 548000 75218 548058 75454
rect 548294 75218 548378 75454
rect 548614 75218 548672 75454
rect 548000 75134 548672 75218
rect 548000 74898 548058 75134
rect 548294 74898 548378 75134
rect 548614 74898 548672 75134
rect 548000 74866 548672 74898
rect 570260 75454 570880 75486
rect 570260 75218 570292 75454
rect 570528 75218 570612 75454
rect 570848 75218 570880 75454
rect 570260 75134 570880 75218
rect 570260 74898 570292 75134
rect 570528 74898 570612 75134
rect 570848 74898 570880 75134
rect 570260 74866 570880 74898
rect 7844 57454 8464 57486
rect 7844 57218 7876 57454
rect 8112 57218 8196 57454
rect 8432 57218 8464 57454
rect 7844 57134 8464 57218
rect 7844 56898 7876 57134
rect 8112 56898 8196 57134
rect 8432 56898 8464 57134
rect 7844 56866 8464 56898
rect 17600 57454 18272 57486
rect 17600 57218 17658 57454
rect 17894 57218 17978 57454
rect 18214 57218 18272 57454
rect 17600 57134 18272 57218
rect 17600 56898 17658 57134
rect 17894 56898 17978 57134
rect 18214 56898 18272 57134
rect 17600 56866 18272 56898
rect 34835 57454 35195 57486
rect 34835 57218 34897 57454
rect 35133 57218 35195 57454
rect 34835 57134 35195 57218
rect 34835 56898 34897 57134
rect 35133 56898 35195 57134
rect 34835 56866 35195 56898
rect 133311 57454 133671 57486
rect 133311 57218 133373 57454
rect 133609 57218 133671 57454
rect 133311 57134 133671 57218
rect 133311 56898 133373 57134
rect 133609 56898 133671 57134
rect 133311 56866 133671 56898
rect 138807 57454 139167 57486
rect 138807 57218 138869 57454
rect 139105 57218 139167 57454
rect 138807 57134 139167 57218
rect 138807 56898 138869 57134
rect 139105 56898 139167 57134
rect 138807 56866 139167 56898
rect 237283 57454 237643 57486
rect 237283 57218 237345 57454
rect 237581 57218 237643 57454
rect 237283 57134 237643 57218
rect 237283 56898 237345 57134
rect 237581 56898 237643 57134
rect 237283 56866 237643 56898
rect 262400 57454 263072 57486
rect 262400 57218 262458 57454
rect 262694 57218 262778 57454
rect 263014 57218 263072 57454
rect 262400 57134 263072 57218
rect 262400 56898 262458 57134
rect 262694 56898 262778 57134
rect 263014 56898 263072 57134
rect 262400 56866 263072 56898
rect 289600 57454 290272 57486
rect 289600 57218 289658 57454
rect 289894 57218 289978 57454
rect 290214 57218 290272 57454
rect 289600 57134 290272 57218
rect 289600 56898 289658 57134
rect 289894 56898 289978 57134
rect 290214 56898 290272 57134
rect 289600 56866 290272 56898
rect 316800 57454 317472 57486
rect 316800 57218 316858 57454
rect 317094 57218 317178 57454
rect 317414 57218 317472 57454
rect 316800 57134 317472 57218
rect 316800 56898 316858 57134
rect 317094 56898 317178 57134
rect 317414 56898 317472 57134
rect 316800 56866 317472 56898
rect 341763 57454 342123 57486
rect 341763 57218 341825 57454
rect 342061 57218 342123 57454
rect 341763 57134 342123 57218
rect 341763 56898 341825 57134
rect 342061 56898 342123 57134
rect 341763 56866 342123 56898
rect 440239 57454 440599 57486
rect 440239 57218 440301 57454
rect 440537 57218 440599 57454
rect 440239 57134 440599 57218
rect 440239 56898 440301 57134
rect 440537 56898 440599 57134
rect 440239 56866 440599 56898
rect 445735 57454 446095 57486
rect 445735 57218 445797 57454
rect 446033 57218 446095 57454
rect 445735 57134 446095 57218
rect 445735 56898 445797 57134
rect 446033 56898 446095 57134
rect 445735 56866 446095 56898
rect 544211 57454 544571 57486
rect 544211 57218 544273 57454
rect 544509 57218 544571 57454
rect 544211 57134 544571 57218
rect 544211 56898 544273 57134
rect 544509 56898 544571 57134
rect 544211 56866 544571 56898
rect 561600 57454 562272 57486
rect 561600 57218 561658 57454
rect 561894 57218 561978 57454
rect 562214 57218 562272 57454
rect 561600 57134 562272 57218
rect 561600 56898 561658 57134
rect 561894 56898 561978 57134
rect 562214 56898 562272 57134
rect 561600 56866 562272 56898
rect 571500 57454 572120 57486
rect 571500 57218 571532 57454
rect 571768 57218 571852 57454
rect 572088 57218 572120 57454
rect 571500 57134 572120 57218
rect 571500 56898 571532 57134
rect 571768 56898 571852 57134
rect 572088 56898 572120 57134
rect 571500 56866 572120 56898
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect 9084 39454 9704 39486
rect 9084 39218 9116 39454
rect 9352 39218 9436 39454
rect 9672 39218 9704 39454
rect 9084 39134 9704 39218
rect 9084 38898 9116 39134
rect 9352 38898 9436 39134
rect 9672 38898 9704 39134
rect 9084 38866 9704 38898
rect 31200 39454 31872 39486
rect 31200 39218 31258 39454
rect 31494 39218 31578 39454
rect 31814 39218 31872 39454
rect 31200 39134 31872 39218
rect 31200 38898 31258 39134
rect 31494 38898 31578 39134
rect 31814 38898 31872 39134
rect 31200 38866 31872 38898
rect 58400 39454 59072 39486
rect 58400 39218 58458 39454
rect 58694 39218 58778 39454
rect 59014 39218 59072 39454
rect 58400 39134 59072 39218
rect 58400 38898 58458 39134
rect 58694 38898 58778 39134
rect 59014 38898 59072 39134
rect 58400 38866 59072 38898
rect 85600 39454 86272 39486
rect 85600 39218 85658 39454
rect 85894 39218 85978 39454
rect 86214 39218 86272 39454
rect 85600 39134 86272 39218
rect 85600 38898 85658 39134
rect 85894 38898 85978 39134
rect 86214 38898 86272 39134
rect 85600 38866 86272 38898
rect 112800 39454 113472 39486
rect 112800 39218 112858 39454
rect 113094 39218 113178 39454
rect 113414 39218 113472 39454
rect 112800 39134 113472 39218
rect 112800 38898 112858 39134
rect 113094 38898 113178 39134
rect 113414 38898 113472 39134
rect 112800 38866 113472 38898
rect 140000 39454 140672 39486
rect 140000 39218 140058 39454
rect 140294 39218 140378 39454
rect 140614 39218 140672 39454
rect 140000 39134 140672 39218
rect 140000 38898 140058 39134
rect 140294 38898 140378 39134
rect 140614 38898 140672 39134
rect 140000 38866 140672 38898
rect 167200 39454 167872 39486
rect 167200 39218 167258 39454
rect 167494 39218 167578 39454
rect 167814 39218 167872 39454
rect 167200 39134 167872 39218
rect 167200 38898 167258 39134
rect 167494 38898 167578 39134
rect 167814 38898 167872 39134
rect 167200 38866 167872 38898
rect 194400 39454 195072 39486
rect 194400 39218 194458 39454
rect 194694 39218 194778 39454
rect 195014 39218 195072 39454
rect 194400 39134 195072 39218
rect 194400 38898 194458 39134
rect 194694 38898 194778 39134
rect 195014 38898 195072 39134
rect 194400 38866 195072 38898
rect 221600 39454 222272 39486
rect 221600 39218 221658 39454
rect 221894 39218 221978 39454
rect 222214 39218 222272 39454
rect 221600 39134 222272 39218
rect 221600 38898 221658 39134
rect 221894 38898 221978 39134
rect 222214 38898 222272 39134
rect 221600 38866 222272 38898
rect 248800 39454 249472 39486
rect 248800 39218 248858 39454
rect 249094 39218 249178 39454
rect 249414 39218 249472 39454
rect 248800 39134 249472 39218
rect 248800 38898 248858 39134
rect 249094 38898 249178 39134
rect 249414 38898 249472 39134
rect 248800 38866 249472 38898
rect 276000 39454 276672 39486
rect 276000 39218 276058 39454
rect 276294 39218 276378 39454
rect 276614 39218 276672 39454
rect 276000 39134 276672 39218
rect 276000 38898 276058 39134
rect 276294 38898 276378 39134
rect 276614 38898 276672 39134
rect 276000 38866 276672 38898
rect 303200 39454 303872 39486
rect 303200 39218 303258 39454
rect 303494 39218 303578 39454
rect 303814 39218 303872 39454
rect 303200 39134 303872 39218
rect 303200 38898 303258 39134
rect 303494 38898 303578 39134
rect 303814 38898 303872 39134
rect 303200 38866 303872 38898
rect 330400 39454 331072 39486
rect 330400 39218 330458 39454
rect 330694 39218 330778 39454
rect 331014 39218 331072 39454
rect 330400 39134 331072 39218
rect 330400 38898 330458 39134
rect 330694 38898 330778 39134
rect 331014 38898 331072 39134
rect 330400 38866 331072 38898
rect 357600 39454 358272 39486
rect 357600 39218 357658 39454
rect 357894 39218 357978 39454
rect 358214 39218 358272 39454
rect 357600 39134 358272 39218
rect 357600 38898 357658 39134
rect 357894 38898 357978 39134
rect 358214 38898 358272 39134
rect 357600 38866 358272 38898
rect 384800 39454 385472 39486
rect 384800 39218 384858 39454
rect 385094 39218 385178 39454
rect 385414 39218 385472 39454
rect 384800 39134 385472 39218
rect 384800 38898 384858 39134
rect 385094 38898 385178 39134
rect 385414 38898 385472 39134
rect 384800 38866 385472 38898
rect 412000 39454 412672 39486
rect 412000 39218 412058 39454
rect 412294 39218 412378 39454
rect 412614 39218 412672 39454
rect 412000 39134 412672 39218
rect 412000 38898 412058 39134
rect 412294 38898 412378 39134
rect 412614 38898 412672 39134
rect 412000 38866 412672 38898
rect 439200 39454 439872 39486
rect 439200 39218 439258 39454
rect 439494 39218 439578 39454
rect 439814 39218 439872 39454
rect 439200 39134 439872 39218
rect 439200 38898 439258 39134
rect 439494 38898 439578 39134
rect 439814 38898 439872 39134
rect 439200 38866 439872 38898
rect 466400 39454 467072 39486
rect 466400 39218 466458 39454
rect 466694 39218 466778 39454
rect 467014 39218 467072 39454
rect 466400 39134 467072 39218
rect 466400 38898 466458 39134
rect 466694 38898 466778 39134
rect 467014 38898 467072 39134
rect 466400 38866 467072 38898
rect 493600 39454 494272 39486
rect 493600 39218 493658 39454
rect 493894 39218 493978 39454
rect 494214 39218 494272 39454
rect 493600 39134 494272 39218
rect 493600 38898 493658 39134
rect 493894 38898 493978 39134
rect 494214 38898 494272 39134
rect 493600 38866 494272 38898
rect 520800 39454 521472 39486
rect 520800 39218 520858 39454
rect 521094 39218 521178 39454
rect 521414 39218 521472 39454
rect 520800 39134 521472 39218
rect 520800 38898 520858 39134
rect 521094 38898 521178 39134
rect 521414 38898 521472 39134
rect 520800 38866 521472 38898
rect 548000 39454 548672 39486
rect 548000 39218 548058 39454
rect 548294 39218 548378 39454
rect 548614 39218 548672 39454
rect 548000 39134 548672 39218
rect 548000 38898 548058 39134
rect 548294 38898 548378 39134
rect 548614 38898 548672 39134
rect 548000 38866 548672 38898
rect 570260 39454 570880 39486
rect 570260 39218 570292 39454
rect 570528 39218 570612 39454
rect 570848 39218 570880 39454
rect 570260 39134 570880 39218
rect 570260 38898 570292 39134
rect 570528 38898 570612 39134
rect 570848 38898 570880 39134
rect 570260 38866 570880 38898
rect 7844 21454 8464 21486
rect 7844 21218 7876 21454
rect 8112 21218 8196 21454
rect 8432 21218 8464 21454
rect 7844 21134 8464 21218
rect 7844 20898 7876 21134
rect 8112 20898 8196 21134
rect 8432 20898 8464 21134
rect 7844 20866 8464 20898
rect 17600 21454 18272 21486
rect 17600 21218 17658 21454
rect 17894 21218 17978 21454
rect 18214 21218 18272 21454
rect 17600 21134 18272 21218
rect 17600 20898 17658 21134
rect 17894 20898 17978 21134
rect 18214 20898 18272 21134
rect 17600 20866 18272 20898
rect 44800 21454 45472 21486
rect 44800 21218 44858 21454
rect 45094 21218 45178 21454
rect 45414 21218 45472 21454
rect 44800 21134 45472 21218
rect 44800 20898 44858 21134
rect 45094 20898 45178 21134
rect 45414 20898 45472 21134
rect 44800 20866 45472 20898
rect 72000 21454 72672 21486
rect 72000 21218 72058 21454
rect 72294 21218 72378 21454
rect 72614 21218 72672 21454
rect 72000 21134 72672 21218
rect 72000 20898 72058 21134
rect 72294 20898 72378 21134
rect 72614 20898 72672 21134
rect 72000 20866 72672 20898
rect 99200 21454 99872 21486
rect 99200 21218 99258 21454
rect 99494 21218 99578 21454
rect 99814 21218 99872 21454
rect 99200 21134 99872 21218
rect 99200 20898 99258 21134
rect 99494 20898 99578 21134
rect 99814 20898 99872 21134
rect 99200 20866 99872 20898
rect 126400 21454 127072 21486
rect 126400 21218 126458 21454
rect 126694 21218 126778 21454
rect 127014 21218 127072 21454
rect 126400 21134 127072 21218
rect 126400 20898 126458 21134
rect 126694 20898 126778 21134
rect 127014 20898 127072 21134
rect 126400 20866 127072 20898
rect 153600 21454 154272 21486
rect 153600 21218 153658 21454
rect 153894 21218 153978 21454
rect 154214 21218 154272 21454
rect 153600 21134 154272 21218
rect 153600 20898 153658 21134
rect 153894 20898 153978 21134
rect 154214 20898 154272 21134
rect 153600 20866 154272 20898
rect 180800 21454 181472 21486
rect 180800 21218 180858 21454
rect 181094 21218 181178 21454
rect 181414 21218 181472 21454
rect 180800 21134 181472 21218
rect 180800 20898 180858 21134
rect 181094 20898 181178 21134
rect 181414 20898 181472 21134
rect 180800 20866 181472 20898
rect 208000 21454 208672 21486
rect 208000 21218 208058 21454
rect 208294 21218 208378 21454
rect 208614 21218 208672 21454
rect 208000 21134 208672 21218
rect 208000 20898 208058 21134
rect 208294 20898 208378 21134
rect 208614 20898 208672 21134
rect 208000 20866 208672 20898
rect 235200 21454 235872 21486
rect 235200 21218 235258 21454
rect 235494 21218 235578 21454
rect 235814 21218 235872 21454
rect 235200 21134 235872 21218
rect 235200 20898 235258 21134
rect 235494 20898 235578 21134
rect 235814 20898 235872 21134
rect 235200 20866 235872 20898
rect 262400 21454 263072 21486
rect 262400 21218 262458 21454
rect 262694 21218 262778 21454
rect 263014 21218 263072 21454
rect 262400 21134 263072 21218
rect 262400 20898 262458 21134
rect 262694 20898 262778 21134
rect 263014 20898 263072 21134
rect 262400 20866 263072 20898
rect 289600 21454 290272 21486
rect 289600 21218 289658 21454
rect 289894 21218 289978 21454
rect 290214 21218 290272 21454
rect 289600 21134 290272 21218
rect 289600 20898 289658 21134
rect 289894 20898 289978 21134
rect 290214 20898 290272 21134
rect 289600 20866 290272 20898
rect 316800 21454 317472 21486
rect 316800 21218 316858 21454
rect 317094 21218 317178 21454
rect 317414 21218 317472 21454
rect 316800 21134 317472 21218
rect 316800 20898 316858 21134
rect 317094 20898 317178 21134
rect 317414 20898 317472 21134
rect 316800 20866 317472 20898
rect 344000 21454 344672 21486
rect 344000 21218 344058 21454
rect 344294 21218 344378 21454
rect 344614 21218 344672 21454
rect 344000 21134 344672 21218
rect 344000 20898 344058 21134
rect 344294 20898 344378 21134
rect 344614 20898 344672 21134
rect 344000 20866 344672 20898
rect 371200 21454 371872 21486
rect 371200 21218 371258 21454
rect 371494 21218 371578 21454
rect 371814 21218 371872 21454
rect 371200 21134 371872 21218
rect 371200 20898 371258 21134
rect 371494 20898 371578 21134
rect 371814 20898 371872 21134
rect 371200 20866 371872 20898
rect 398400 21454 399072 21486
rect 398400 21218 398458 21454
rect 398694 21218 398778 21454
rect 399014 21218 399072 21454
rect 398400 21134 399072 21218
rect 398400 20898 398458 21134
rect 398694 20898 398778 21134
rect 399014 20898 399072 21134
rect 398400 20866 399072 20898
rect 425600 21454 426272 21486
rect 425600 21218 425658 21454
rect 425894 21218 425978 21454
rect 426214 21218 426272 21454
rect 425600 21134 426272 21218
rect 425600 20898 425658 21134
rect 425894 20898 425978 21134
rect 426214 20898 426272 21134
rect 425600 20866 426272 20898
rect 452800 21454 453472 21486
rect 452800 21218 452858 21454
rect 453094 21218 453178 21454
rect 453414 21218 453472 21454
rect 452800 21134 453472 21218
rect 452800 20898 452858 21134
rect 453094 20898 453178 21134
rect 453414 20898 453472 21134
rect 452800 20866 453472 20898
rect 480000 21454 480672 21486
rect 480000 21218 480058 21454
rect 480294 21218 480378 21454
rect 480614 21218 480672 21454
rect 480000 21134 480672 21218
rect 480000 20898 480058 21134
rect 480294 20898 480378 21134
rect 480614 20898 480672 21134
rect 480000 20866 480672 20898
rect 507200 21454 507872 21486
rect 507200 21218 507258 21454
rect 507494 21218 507578 21454
rect 507814 21218 507872 21454
rect 507200 21134 507872 21218
rect 507200 20898 507258 21134
rect 507494 20898 507578 21134
rect 507814 20898 507872 21134
rect 507200 20866 507872 20898
rect 534400 21454 535072 21486
rect 534400 21218 534458 21454
rect 534694 21218 534778 21454
rect 535014 21218 535072 21454
rect 534400 21134 535072 21218
rect 534400 20898 534458 21134
rect 534694 20898 534778 21134
rect 535014 20898 535072 21134
rect 534400 20866 535072 20898
rect 561600 21454 562272 21486
rect 561600 21218 561658 21454
rect 561894 21218 561978 21454
rect 562214 21218 562272 21454
rect 561600 21134 562272 21218
rect 561600 20898 561658 21134
rect 561894 20898 561978 21134
rect 562214 20898 562272 21134
rect 561600 20866 562272 20898
rect 571500 21454 572120 21486
rect 571500 21218 571532 21454
rect 571768 21218 571852 21454
rect 572088 21218 572120 21454
rect 571500 21134 572120 21218
rect 571500 20898 571532 21134
rect 571768 20898 571852 21134
rect 572088 20898 572120 21134
rect 571500 20866 572120 20898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 -346 2414 2000
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 2000
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 2000
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 2000
rect 19794 -1306 20414 2000
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 -3226 24134 2000
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 -5146 27854 2000
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 2000
rect 37794 -346 38414 2000
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 -2266 42134 2000
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 -4186 45854 2000
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 2000
rect 55794 -1306 56414 2000
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 -3226 60134 2000
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 -5146 63854 2000
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 2000
rect 73794 -346 74414 2000
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 -2266 78134 2000
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 -4186 81854 2000
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 2000
rect 91794 -1306 92414 2000
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 -3226 96134 2000
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 -5146 99854 2000
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 2000
rect 109794 -346 110414 2000
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 -2266 114134 2000
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 -4186 117854 2000
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 2000
rect 127794 -1306 128414 2000
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 -3226 132134 2000
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 -5146 135854 2000
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 2000
rect 145794 -346 146414 2000
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 -2266 150134 2000
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 -4186 153854 2000
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 2000
rect 163794 -1306 164414 2000
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 -3226 168134 2000
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 -5146 171854 2000
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 2000
rect 181794 -346 182414 2000
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 -2266 186134 2000
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 -4186 189854 2000
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 2000
rect 199794 -1306 200414 2000
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 -3226 204134 2000
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 -5146 207854 2000
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 2000
rect 217794 -346 218414 2000
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 -2266 222134 2000
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 -4186 225854 2000
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 2000
rect 235794 -1306 236414 2000
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 -3226 240134 2000
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 -5146 243854 2000
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 2000
rect 253794 -346 254414 2000
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 -2266 258134 2000
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 -4186 261854 2000
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 2000
rect 271794 -1306 272414 2000
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 -3226 276134 2000
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 -5146 279854 2000
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 2000
rect 289794 -346 290414 2000
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 -2266 294134 2000
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 -4186 297854 2000
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 2000
rect 307794 -1306 308414 2000
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 -3226 312134 2000
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 -5146 315854 2000
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 2000
rect 325794 -346 326414 2000
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 -2266 330134 2000
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 -4186 333854 2000
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 2000
rect 343794 -1306 344414 2000
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 -3226 348134 2000
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 -5146 351854 2000
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 2000
rect 361794 -346 362414 2000
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 -2266 366134 2000
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 -4186 369854 2000
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 2000
rect 379794 -1306 380414 2000
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 -3226 384134 2000
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 -5146 387854 2000
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 2000
rect 397794 -346 398414 2000
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 -2266 402134 2000
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 -4186 405854 2000
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 2000
rect 415794 -1306 416414 2000
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 -3226 420134 2000
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 -5146 423854 2000
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 2000
rect 433794 -346 434414 2000
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 -2266 438134 2000
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 -4186 441854 2000
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 2000
rect 451794 -1306 452414 2000
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 -3226 456134 2000
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 -5146 459854 2000
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 2000
rect 469794 -346 470414 2000
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 -2266 474134 2000
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 -4186 477854 2000
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 2000
rect 487794 -1306 488414 2000
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 -3226 492134 2000
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 -5146 495854 2000
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 2000
rect 505794 -346 506414 2000
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 -2266 510134 2000
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 -4186 513854 2000
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 2000
rect 523794 -1306 524414 2000
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 -3226 528134 2000
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 -5146 531854 2000
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 2000
rect 541794 -346 542414 2000
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 -2266 546134 2000
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 -4186 549854 2000
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 2000
rect 559794 -1306 560414 2000
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 -3226 564134 2000
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 -5146 567854 2000
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 2000
rect 577794 -346 578414 2000
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect 9116 687218 9352 687454
rect 9436 687218 9672 687454
rect 9116 686898 9352 687134
rect 9436 686898 9672 687134
rect 31258 687218 31494 687454
rect 31578 687218 31814 687454
rect 31258 686898 31494 687134
rect 31578 686898 31814 687134
rect 58458 687218 58694 687454
rect 58778 687218 59014 687454
rect 58458 686898 58694 687134
rect 58778 686898 59014 687134
rect 85658 687218 85894 687454
rect 85978 687218 86214 687454
rect 85658 686898 85894 687134
rect 85978 686898 86214 687134
rect 112858 687218 113094 687454
rect 113178 687218 113414 687454
rect 112858 686898 113094 687134
rect 113178 686898 113414 687134
rect 140058 687218 140294 687454
rect 140378 687218 140614 687454
rect 140058 686898 140294 687134
rect 140378 686898 140614 687134
rect 167258 687218 167494 687454
rect 167578 687218 167814 687454
rect 167258 686898 167494 687134
rect 167578 686898 167814 687134
rect 194458 687218 194694 687454
rect 194778 687218 195014 687454
rect 194458 686898 194694 687134
rect 194778 686898 195014 687134
rect 221658 687218 221894 687454
rect 221978 687218 222214 687454
rect 221658 686898 221894 687134
rect 221978 686898 222214 687134
rect 248858 687218 249094 687454
rect 249178 687218 249414 687454
rect 248858 686898 249094 687134
rect 249178 686898 249414 687134
rect 276058 687218 276294 687454
rect 276378 687218 276614 687454
rect 276058 686898 276294 687134
rect 276378 686898 276614 687134
rect 303258 687218 303494 687454
rect 303578 687218 303814 687454
rect 303258 686898 303494 687134
rect 303578 686898 303814 687134
rect 330458 687218 330694 687454
rect 330778 687218 331014 687454
rect 330458 686898 330694 687134
rect 330778 686898 331014 687134
rect 357658 687218 357894 687454
rect 357978 687218 358214 687454
rect 357658 686898 357894 687134
rect 357978 686898 358214 687134
rect 384858 687218 385094 687454
rect 385178 687218 385414 687454
rect 384858 686898 385094 687134
rect 385178 686898 385414 687134
rect 412058 687218 412294 687454
rect 412378 687218 412614 687454
rect 412058 686898 412294 687134
rect 412378 686898 412614 687134
rect 439258 687218 439494 687454
rect 439578 687218 439814 687454
rect 439258 686898 439494 687134
rect 439578 686898 439814 687134
rect 466458 687218 466694 687454
rect 466778 687218 467014 687454
rect 466458 686898 466694 687134
rect 466778 686898 467014 687134
rect 493658 687218 493894 687454
rect 493978 687218 494214 687454
rect 493658 686898 493894 687134
rect 493978 686898 494214 687134
rect 520858 687218 521094 687454
rect 521178 687218 521414 687454
rect 520858 686898 521094 687134
rect 521178 686898 521414 687134
rect 548058 687218 548294 687454
rect 548378 687218 548614 687454
rect 548058 686898 548294 687134
rect 548378 686898 548614 687134
rect 570292 687218 570528 687454
rect 570612 687218 570848 687454
rect 570292 686898 570528 687134
rect 570612 686898 570848 687134
rect 7876 669218 8112 669454
rect 8196 669218 8432 669454
rect 7876 668898 8112 669134
rect 8196 668898 8432 669134
rect 17658 669218 17894 669454
rect 17978 669218 18214 669454
rect 17658 668898 17894 669134
rect 17978 668898 18214 669134
rect 44858 669218 45094 669454
rect 45178 669218 45414 669454
rect 44858 668898 45094 669134
rect 45178 668898 45414 669134
rect 72058 669218 72294 669454
rect 72378 669218 72614 669454
rect 72058 668898 72294 669134
rect 72378 668898 72614 669134
rect 99258 669218 99494 669454
rect 99578 669218 99814 669454
rect 99258 668898 99494 669134
rect 99578 668898 99814 669134
rect 126458 669218 126694 669454
rect 126778 669218 127014 669454
rect 126458 668898 126694 669134
rect 126778 668898 127014 669134
rect 153658 669218 153894 669454
rect 153978 669218 154214 669454
rect 153658 668898 153894 669134
rect 153978 668898 154214 669134
rect 180858 669218 181094 669454
rect 181178 669218 181414 669454
rect 180858 668898 181094 669134
rect 181178 668898 181414 669134
rect 208058 669218 208294 669454
rect 208378 669218 208614 669454
rect 208058 668898 208294 669134
rect 208378 668898 208614 669134
rect 235258 669218 235494 669454
rect 235578 669218 235814 669454
rect 235258 668898 235494 669134
rect 235578 668898 235814 669134
rect 262458 669218 262694 669454
rect 262778 669218 263014 669454
rect 262458 668898 262694 669134
rect 262778 668898 263014 669134
rect 289658 669218 289894 669454
rect 289978 669218 290214 669454
rect 289658 668898 289894 669134
rect 289978 668898 290214 669134
rect 316858 669218 317094 669454
rect 317178 669218 317414 669454
rect 316858 668898 317094 669134
rect 317178 668898 317414 669134
rect 344058 669218 344294 669454
rect 344378 669218 344614 669454
rect 344058 668898 344294 669134
rect 344378 668898 344614 669134
rect 371258 669218 371494 669454
rect 371578 669218 371814 669454
rect 371258 668898 371494 669134
rect 371578 668898 371814 669134
rect 398458 669218 398694 669454
rect 398778 669218 399014 669454
rect 398458 668898 398694 669134
rect 398778 668898 399014 669134
rect 425658 669218 425894 669454
rect 425978 669218 426214 669454
rect 425658 668898 425894 669134
rect 425978 668898 426214 669134
rect 452858 669218 453094 669454
rect 453178 669218 453414 669454
rect 452858 668898 453094 669134
rect 453178 668898 453414 669134
rect 480058 669218 480294 669454
rect 480378 669218 480614 669454
rect 480058 668898 480294 669134
rect 480378 668898 480614 669134
rect 507258 669218 507494 669454
rect 507578 669218 507814 669454
rect 507258 668898 507494 669134
rect 507578 668898 507814 669134
rect 534458 669218 534694 669454
rect 534778 669218 535014 669454
rect 534458 668898 534694 669134
rect 534778 668898 535014 669134
rect 561658 669218 561894 669454
rect 561978 669218 562214 669454
rect 561658 668898 561894 669134
rect 561978 668898 562214 669134
rect 571532 669218 571768 669454
rect 571852 669218 572088 669454
rect 571532 668898 571768 669134
rect 571852 668898 572088 669134
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect 9116 651218 9352 651454
rect 9436 651218 9672 651454
rect 9116 650898 9352 651134
rect 9436 650898 9672 651134
rect 31258 651218 31494 651454
rect 31578 651218 31814 651454
rect 31258 650898 31494 651134
rect 31578 650898 31814 651134
rect 58458 651218 58694 651454
rect 58778 651218 59014 651454
rect 58458 650898 58694 651134
rect 58778 650898 59014 651134
rect 85658 651218 85894 651454
rect 85978 651218 86214 651454
rect 85658 650898 85894 651134
rect 85978 650898 86214 651134
rect 112858 651218 113094 651454
rect 113178 651218 113414 651454
rect 112858 650898 113094 651134
rect 113178 650898 113414 651134
rect 140058 651218 140294 651454
rect 140378 651218 140614 651454
rect 140058 650898 140294 651134
rect 140378 650898 140614 651134
rect 167258 651218 167494 651454
rect 167578 651218 167814 651454
rect 167258 650898 167494 651134
rect 167578 650898 167814 651134
rect 194458 651218 194694 651454
rect 194778 651218 195014 651454
rect 194458 650898 194694 651134
rect 194778 650898 195014 651134
rect 221658 651218 221894 651454
rect 221978 651218 222214 651454
rect 221658 650898 221894 651134
rect 221978 650898 222214 651134
rect 248858 651218 249094 651454
rect 249178 651218 249414 651454
rect 248858 650898 249094 651134
rect 249178 650898 249414 651134
rect 276058 651218 276294 651454
rect 276378 651218 276614 651454
rect 276058 650898 276294 651134
rect 276378 650898 276614 651134
rect 303258 651218 303494 651454
rect 303578 651218 303814 651454
rect 303258 650898 303494 651134
rect 303578 650898 303814 651134
rect 330458 651218 330694 651454
rect 330778 651218 331014 651454
rect 330458 650898 330694 651134
rect 330778 650898 331014 651134
rect 357658 651218 357894 651454
rect 357978 651218 358214 651454
rect 357658 650898 357894 651134
rect 357978 650898 358214 651134
rect 384858 651218 385094 651454
rect 385178 651218 385414 651454
rect 384858 650898 385094 651134
rect 385178 650898 385414 651134
rect 412058 651218 412294 651454
rect 412378 651218 412614 651454
rect 412058 650898 412294 651134
rect 412378 650898 412614 651134
rect 439258 651218 439494 651454
rect 439578 651218 439814 651454
rect 439258 650898 439494 651134
rect 439578 650898 439814 651134
rect 466458 651218 466694 651454
rect 466778 651218 467014 651454
rect 466458 650898 466694 651134
rect 466778 650898 467014 651134
rect 493658 651218 493894 651454
rect 493978 651218 494214 651454
rect 493658 650898 493894 651134
rect 493978 650898 494214 651134
rect 520858 651218 521094 651454
rect 521178 651218 521414 651454
rect 520858 650898 521094 651134
rect 521178 650898 521414 651134
rect 548058 651218 548294 651454
rect 548378 651218 548614 651454
rect 548058 650898 548294 651134
rect 548378 650898 548614 651134
rect 570292 651218 570528 651454
rect 570612 651218 570848 651454
rect 570292 650898 570528 651134
rect 570612 650898 570848 651134
rect 7876 633218 8112 633454
rect 8196 633218 8432 633454
rect 7876 632898 8112 633134
rect 8196 632898 8432 633134
rect 17658 633218 17894 633454
rect 17978 633218 18214 633454
rect 17658 632898 17894 633134
rect 17978 632898 18214 633134
rect 44858 633218 45094 633454
rect 45178 633218 45414 633454
rect 44858 632898 45094 633134
rect 45178 632898 45414 633134
rect 72058 633218 72294 633454
rect 72378 633218 72614 633454
rect 72058 632898 72294 633134
rect 72378 632898 72614 633134
rect 99258 633218 99494 633454
rect 99578 633218 99814 633454
rect 99258 632898 99494 633134
rect 99578 632898 99814 633134
rect 126458 633218 126694 633454
rect 126778 633218 127014 633454
rect 126458 632898 126694 633134
rect 126778 632898 127014 633134
rect 153658 633218 153894 633454
rect 153978 633218 154214 633454
rect 153658 632898 153894 633134
rect 153978 632898 154214 633134
rect 180858 633218 181094 633454
rect 181178 633218 181414 633454
rect 180858 632898 181094 633134
rect 181178 632898 181414 633134
rect 208058 633218 208294 633454
rect 208378 633218 208614 633454
rect 208058 632898 208294 633134
rect 208378 632898 208614 633134
rect 235258 633218 235494 633454
rect 235578 633218 235814 633454
rect 235258 632898 235494 633134
rect 235578 632898 235814 633134
rect 262458 633218 262694 633454
rect 262778 633218 263014 633454
rect 262458 632898 262694 633134
rect 262778 632898 263014 633134
rect 289658 633218 289894 633454
rect 289978 633218 290214 633454
rect 289658 632898 289894 633134
rect 289978 632898 290214 633134
rect 316858 633218 317094 633454
rect 317178 633218 317414 633454
rect 316858 632898 317094 633134
rect 317178 632898 317414 633134
rect 344058 633218 344294 633454
rect 344378 633218 344614 633454
rect 344058 632898 344294 633134
rect 344378 632898 344614 633134
rect 371258 633218 371494 633454
rect 371578 633218 371814 633454
rect 371258 632898 371494 633134
rect 371578 632898 371814 633134
rect 398458 633218 398694 633454
rect 398778 633218 399014 633454
rect 398458 632898 398694 633134
rect 398778 632898 399014 633134
rect 425658 633218 425894 633454
rect 425978 633218 426214 633454
rect 425658 632898 425894 633134
rect 425978 632898 426214 633134
rect 452858 633218 453094 633454
rect 453178 633218 453414 633454
rect 452858 632898 453094 633134
rect 453178 632898 453414 633134
rect 480058 633218 480294 633454
rect 480378 633218 480614 633454
rect 480058 632898 480294 633134
rect 480378 632898 480614 633134
rect 507258 633218 507494 633454
rect 507578 633218 507814 633454
rect 507258 632898 507494 633134
rect 507578 632898 507814 633134
rect 534458 633218 534694 633454
rect 534778 633218 535014 633454
rect 534458 632898 534694 633134
rect 534778 632898 535014 633134
rect 561658 633218 561894 633454
rect 561978 633218 562214 633454
rect 561658 632898 561894 633134
rect 561978 632898 562214 633134
rect 571532 633218 571768 633454
rect 571852 633218 572088 633454
rect 571532 632898 571768 633134
rect 571852 632898 572088 633134
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect 9116 615218 9352 615454
rect 9436 615218 9672 615454
rect 9116 614898 9352 615134
rect 9436 614898 9672 615134
rect 31258 615218 31494 615454
rect 31578 615218 31814 615454
rect 31258 614898 31494 615134
rect 31578 614898 31814 615134
rect 58458 615218 58694 615454
rect 58778 615218 59014 615454
rect 58458 614898 58694 615134
rect 58778 614898 59014 615134
rect 85658 615218 85894 615454
rect 85978 615218 86214 615454
rect 85658 614898 85894 615134
rect 85978 614898 86214 615134
rect 112858 615218 113094 615454
rect 113178 615218 113414 615454
rect 112858 614898 113094 615134
rect 113178 614898 113414 615134
rect 140058 615218 140294 615454
rect 140378 615218 140614 615454
rect 140058 614898 140294 615134
rect 140378 614898 140614 615134
rect 167258 615218 167494 615454
rect 167578 615218 167814 615454
rect 167258 614898 167494 615134
rect 167578 614898 167814 615134
rect 194458 615218 194694 615454
rect 194778 615218 195014 615454
rect 194458 614898 194694 615134
rect 194778 614898 195014 615134
rect 221658 615218 221894 615454
rect 221978 615218 222214 615454
rect 221658 614898 221894 615134
rect 221978 614898 222214 615134
rect 248858 615218 249094 615454
rect 249178 615218 249414 615454
rect 248858 614898 249094 615134
rect 249178 614898 249414 615134
rect 276058 615218 276294 615454
rect 276378 615218 276614 615454
rect 276058 614898 276294 615134
rect 276378 614898 276614 615134
rect 303258 615218 303494 615454
rect 303578 615218 303814 615454
rect 303258 614898 303494 615134
rect 303578 614898 303814 615134
rect 330458 615218 330694 615454
rect 330778 615218 331014 615454
rect 330458 614898 330694 615134
rect 330778 614898 331014 615134
rect 357658 615218 357894 615454
rect 357978 615218 358214 615454
rect 357658 614898 357894 615134
rect 357978 614898 358214 615134
rect 384858 615218 385094 615454
rect 385178 615218 385414 615454
rect 384858 614898 385094 615134
rect 385178 614898 385414 615134
rect 412058 615218 412294 615454
rect 412378 615218 412614 615454
rect 412058 614898 412294 615134
rect 412378 614898 412614 615134
rect 439258 615218 439494 615454
rect 439578 615218 439814 615454
rect 439258 614898 439494 615134
rect 439578 614898 439814 615134
rect 466458 615218 466694 615454
rect 466778 615218 467014 615454
rect 466458 614898 466694 615134
rect 466778 614898 467014 615134
rect 493658 615218 493894 615454
rect 493978 615218 494214 615454
rect 493658 614898 493894 615134
rect 493978 614898 494214 615134
rect 520858 615218 521094 615454
rect 521178 615218 521414 615454
rect 520858 614898 521094 615134
rect 521178 614898 521414 615134
rect 548058 615218 548294 615454
rect 548378 615218 548614 615454
rect 548058 614898 548294 615134
rect 548378 614898 548614 615134
rect 570292 615218 570528 615454
rect 570612 615218 570848 615454
rect 570292 614898 570528 615134
rect 570612 614898 570848 615134
rect 7876 597218 8112 597454
rect 8196 597218 8432 597454
rect 7876 596898 8112 597134
rect 8196 596898 8432 597134
rect 17658 597218 17894 597454
rect 17978 597218 18214 597454
rect 17658 596898 17894 597134
rect 17978 596898 18214 597134
rect 34897 597218 35133 597454
rect 34897 596898 35133 597134
rect 133373 597218 133609 597454
rect 133373 596898 133609 597134
rect 138869 597218 139105 597454
rect 138869 596898 139105 597134
rect 237345 597218 237581 597454
rect 237345 596898 237581 597134
rect 262458 597218 262694 597454
rect 262778 597218 263014 597454
rect 262458 596898 262694 597134
rect 262778 596898 263014 597134
rect 289658 597218 289894 597454
rect 289978 597218 290214 597454
rect 289658 596898 289894 597134
rect 289978 596898 290214 597134
rect 316858 597218 317094 597454
rect 317178 597218 317414 597454
rect 316858 596898 317094 597134
rect 317178 596898 317414 597134
rect 341825 597218 342061 597454
rect 341825 596898 342061 597134
rect 440301 597218 440537 597454
rect 440301 596898 440537 597134
rect 445797 597218 446033 597454
rect 445797 596898 446033 597134
rect 544273 597218 544509 597454
rect 544273 596898 544509 597134
rect 561658 597218 561894 597454
rect 561978 597218 562214 597454
rect 561658 596898 561894 597134
rect 561978 596898 562214 597134
rect 571532 597218 571768 597454
rect 571852 597218 572088 597454
rect 571532 596898 571768 597134
rect 571852 596898 572088 597134
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect 9116 579218 9352 579454
rect 9436 579218 9672 579454
rect 9116 578898 9352 579134
rect 9436 578898 9672 579134
rect 31258 579218 31494 579454
rect 31578 579218 31814 579454
rect 31258 578898 31494 579134
rect 31578 578898 31814 579134
rect 35617 579218 35853 579454
rect 35617 578898 35853 579134
rect 132653 579218 132889 579454
rect 132653 578898 132889 579134
rect 139589 579218 139825 579454
rect 139589 578898 139825 579134
rect 236625 579218 236861 579454
rect 236625 578898 236861 579134
rect 248858 579218 249094 579454
rect 249178 579218 249414 579454
rect 248858 578898 249094 579134
rect 249178 578898 249414 579134
rect 276058 579218 276294 579454
rect 276378 579218 276614 579454
rect 276058 578898 276294 579134
rect 276378 578898 276614 579134
rect 303258 579218 303494 579454
rect 303578 579218 303814 579454
rect 303258 578898 303494 579134
rect 303578 578898 303814 579134
rect 330458 579218 330694 579454
rect 330778 579218 331014 579454
rect 330458 578898 330694 579134
rect 330778 578898 331014 579134
rect 342545 579218 342781 579454
rect 342545 578898 342781 579134
rect 439581 579218 439817 579454
rect 439581 578898 439817 579134
rect 446517 579218 446753 579454
rect 446517 578898 446753 579134
rect 543553 579218 543789 579454
rect 543553 578898 543789 579134
rect 548058 579218 548294 579454
rect 548378 579218 548614 579454
rect 548058 578898 548294 579134
rect 548378 578898 548614 579134
rect 570292 579218 570528 579454
rect 570612 579218 570848 579454
rect 570292 578898 570528 579134
rect 570612 578898 570848 579134
rect 7876 561218 8112 561454
rect 8196 561218 8432 561454
rect 7876 560898 8112 561134
rect 8196 560898 8432 561134
rect 17658 561218 17894 561454
rect 17978 561218 18214 561454
rect 17658 560898 17894 561134
rect 17978 560898 18214 561134
rect 34897 561218 35133 561454
rect 34897 560898 35133 561134
rect 133373 561218 133609 561454
rect 133373 560898 133609 561134
rect 138869 561218 139105 561454
rect 138869 560898 139105 561134
rect 237345 561218 237581 561454
rect 237345 560898 237581 561134
rect 262458 561218 262694 561454
rect 262778 561218 263014 561454
rect 262458 560898 262694 561134
rect 262778 560898 263014 561134
rect 289658 561218 289894 561454
rect 289978 561218 290214 561454
rect 289658 560898 289894 561134
rect 289978 560898 290214 561134
rect 316858 561218 317094 561454
rect 317178 561218 317414 561454
rect 316858 560898 317094 561134
rect 317178 560898 317414 561134
rect 341825 561218 342061 561454
rect 341825 560898 342061 561134
rect 440301 561218 440537 561454
rect 440301 560898 440537 561134
rect 445797 561218 446033 561454
rect 445797 560898 446033 561134
rect 544273 561218 544509 561454
rect 544273 560898 544509 561134
rect 561658 561218 561894 561454
rect 561978 561218 562214 561454
rect 561658 560898 561894 561134
rect 561978 560898 562214 561134
rect 571532 561218 571768 561454
rect 571852 561218 572088 561454
rect 571532 560898 571768 561134
rect 571852 560898 572088 561134
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect 9116 543218 9352 543454
rect 9436 543218 9672 543454
rect 9116 542898 9352 543134
rect 9436 542898 9672 543134
rect 31258 543218 31494 543454
rect 31578 543218 31814 543454
rect 31258 542898 31494 543134
rect 31578 542898 31814 543134
rect 35617 543218 35853 543454
rect 35617 542898 35853 543134
rect 132653 543218 132889 543454
rect 132653 542898 132889 543134
rect 139589 543218 139825 543454
rect 139589 542898 139825 543134
rect 236625 543218 236861 543454
rect 236625 542898 236861 543134
rect 248858 543218 249094 543454
rect 249178 543218 249414 543454
rect 248858 542898 249094 543134
rect 249178 542898 249414 543134
rect 276058 543218 276294 543454
rect 276378 543218 276614 543454
rect 276058 542898 276294 543134
rect 276378 542898 276614 543134
rect 303258 543218 303494 543454
rect 303578 543218 303814 543454
rect 303258 542898 303494 543134
rect 303578 542898 303814 543134
rect 330458 543218 330694 543454
rect 330778 543218 331014 543454
rect 330458 542898 330694 543134
rect 330778 542898 331014 543134
rect 342545 543218 342781 543454
rect 342545 542898 342781 543134
rect 439581 543218 439817 543454
rect 439581 542898 439817 543134
rect 446517 543218 446753 543454
rect 446517 542898 446753 543134
rect 543553 543218 543789 543454
rect 543553 542898 543789 543134
rect 548058 543218 548294 543454
rect 548378 543218 548614 543454
rect 548058 542898 548294 543134
rect 548378 542898 548614 543134
rect 570292 543218 570528 543454
rect 570612 543218 570848 543454
rect 570292 542898 570528 543134
rect 570612 542898 570848 543134
rect 7876 525218 8112 525454
rect 8196 525218 8432 525454
rect 7876 524898 8112 525134
rect 8196 524898 8432 525134
rect 17658 525218 17894 525454
rect 17978 525218 18214 525454
rect 17658 524898 17894 525134
rect 17978 524898 18214 525134
rect 44858 525218 45094 525454
rect 45178 525218 45414 525454
rect 44858 524898 45094 525134
rect 45178 524898 45414 525134
rect 72058 525218 72294 525454
rect 72378 525218 72614 525454
rect 72058 524898 72294 525134
rect 72378 524898 72614 525134
rect 99258 525218 99494 525454
rect 99578 525218 99814 525454
rect 99258 524898 99494 525134
rect 99578 524898 99814 525134
rect 126458 525218 126694 525454
rect 126778 525218 127014 525454
rect 126458 524898 126694 525134
rect 126778 524898 127014 525134
rect 153658 525218 153894 525454
rect 153978 525218 154214 525454
rect 153658 524898 153894 525134
rect 153978 524898 154214 525134
rect 180858 525218 181094 525454
rect 181178 525218 181414 525454
rect 180858 524898 181094 525134
rect 181178 524898 181414 525134
rect 208058 525218 208294 525454
rect 208378 525218 208614 525454
rect 208058 524898 208294 525134
rect 208378 524898 208614 525134
rect 235258 525218 235494 525454
rect 235578 525218 235814 525454
rect 235258 524898 235494 525134
rect 235578 524898 235814 525134
rect 262458 525218 262694 525454
rect 262778 525218 263014 525454
rect 262458 524898 262694 525134
rect 262778 524898 263014 525134
rect 289658 525218 289894 525454
rect 289978 525218 290214 525454
rect 289658 524898 289894 525134
rect 289978 524898 290214 525134
rect 316858 525218 317094 525454
rect 317178 525218 317414 525454
rect 316858 524898 317094 525134
rect 317178 524898 317414 525134
rect 344058 525218 344294 525454
rect 344378 525218 344614 525454
rect 344058 524898 344294 525134
rect 344378 524898 344614 525134
rect 371258 525218 371494 525454
rect 371578 525218 371814 525454
rect 371258 524898 371494 525134
rect 371578 524898 371814 525134
rect 398458 525218 398694 525454
rect 398778 525218 399014 525454
rect 398458 524898 398694 525134
rect 398778 524898 399014 525134
rect 425658 525218 425894 525454
rect 425978 525218 426214 525454
rect 425658 524898 425894 525134
rect 425978 524898 426214 525134
rect 452858 525218 453094 525454
rect 453178 525218 453414 525454
rect 452858 524898 453094 525134
rect 453178 524898 453414 525134
rect 480058 525218 480294 525454
rect 480378 525218 480614 525454
rect 480058 524898 480294 525134
rect 480378 524898 480614 525134
rect 507258 525218 507494 525454
rect 507578 525218 507814 525454
rect 507258 524898 507494 525134
rect 507578 524898 507814 525134
rect 534458 525218 534694 525454
rect 534778 525218 535014 525454
rect 534458 524898 534694 525134
rect 534778 524898 535014 525134
rect 561658 525218 561894 525454
rect 561978 525218 562214 525454
rect 561658 524898 561894 525134
rect 561978 524898 562214 525134
rect 571532 525218 571768 525454
rect 571852 525218 572088 525454
rect 571532 524898 571768 525134
rect 571852 524898 572088 525134
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect 9116 507218 9352 507454
rect 9436 507218 9672 507454
rect 9116 506898 9352 507134
rect 9436 506898 9672 507134
rect 31258 507218 31494 507454
rect 31578 507218 31814 507454
rect 31258 506898 31494 507134
rect 31578 506898 31814 507134
rect 35617 507218 35853 507454
rect 35617 506898 35853 507134
rect 132653 507218 132889 507454
rect 132653 506898 132889 507134
rect 139589 507218 139825 507454
rect 139589 506898 139825 507134
rect 236625 507218 236861 507454
rect 236625 506898 236861 507134
rect 248858 507218 249094 507454
rect 249178 507218 249414 507454
rect 248858 506898 249094 507134
rect 249178 506898 249414 507134
rect 276058 507218 276294 507454
rect 276378 507218 276614 507454
rect 276058 506898 276294 507134
rect 276378 506898 276614 507134
rect 303258 507218 303494 507454
rect 303578 507218 303814 507454
rect 303258 506898 303494 507134
rect 303578 506898 303814 507134
rect 330458 507218 330694 507454
rect 330778 507218 331014 507454
rect 330458 506898 330694 507134
rect 330778 506898 331014 507134
rect 342545 507218 342781 507454
rect 342545 506898 342781 507134
rect 439581 507218 439817 507454
rect 439581 506898 439817 507134
rect 446517 507218 446753 507454
rect 446517 506898 446753 507134
rect 543553 507218 543789 507454
rect 543553 506898 543789 507134
rect 548058 507218 548294 507454
rect 548378 507218 548614 507454
rect 548058 506898 548294 507134
rect 548378 506898 548614 507134
rect 570292 507218 570528 507454
rect 570612 507218 570848 507454
rect 570292 506898 570528 507134
rect 570612 506898 570848 507134
rect 7876 489218 8112 489454
rect 8196 489218 8432 489454
rect 7876 488898 8112 489134
rect 8196 488898 8432 489134
rect 17658 489218 17894 489454
rect 17978 489218 18214 489454
rect 17658 488898 17894 489134
rect 17978 488898 18214 489134
rect 34897 489218 35133 489454
rect 34897 488898 35133 489134
rect 133373 489218 133609 489454
rect 133373 488898 133609 489134
rect 138869 489218 139105 489454
rect 138869 488898 139105 489134
rect 237345 489218 237581 489454
rect 237345 488898 237581 489134
rect 262458 489218 262694 489454
rect 262778 489218 263014 489454
rect 262458 488898 262694 489134
rect 262778 488898 263014 489134
rect 289658 489218 289894 489454
rect 289978 489218 290214 489454
rect 289658 488898 289894 489134
rect 289978 488898 290214 489134
rect 316858 489218 317094 489454
rect 317178 489218 317414 489454
rect 316858 488898 317094 489134
rect 317178 488898 317414 489134
rect 341825 489218 342061 489454
rect 341825 488898 342061 489134
rect 440301 489218 440537 489454
rect 440301 488898 440537 489134
rect 445797 489218 446033 489454
rect 445797 488898 446033 489134
rect 544273 489218 544509 489454
rect 544273 488898 544509 489134
rect 561658 489218 561894 489454
rect 561978 489218 562214 489454
rect 561658 488898 561894 489134
rect 561978 488898 562214 489134
rect 571532 489218 571768 489454
rect 571852 489218 572088 489454
rect 571532 488898 571768 489134
rect 571852 488898 572088 489134
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect 9116 471218 9352 471454
rect 9436 471218 9672 471454
rect 9116 470898 9352 471134
rect 9436 470898 9672 471134
rect 31258 471218 31494 471454
rect 31578 471218 31814 471454
rect 31258 470898 31494 471134
rect 31578 470898 31814 471134
rect 35617 471218 35853 471454
rect 35617 470898 35853 471134
rect 132653 471218 132889 471454
rect 132653 470898 132889 471134
rect 139589 471218 139825 471454
rect 139589 470898 139825 471134
rect 236625 471218 236861 471454
rect 236625 470898 236861 471134
rect 248858 471218 249094 471454
rect 249178 471218 249414 471454
rect 248858 470898 249094 471134
rect 249178 470898 249414 471134
rect 276058 471218 276294 471454
rect 276378 471218 276614 471454
rect 276058 470898 276294 471134
rect 276378 470898 276614 471134
rect 303258 471218 303494 471454
rect 303578 471218 303814 471454
rect 303258 470898 303494 471134
rect 303578 470898 303814 471134
rect 330458 471218 330694 471454
rect 330778 471218 331014 471454
rect 330458 470898 330694 471134
rect 330778 470898 331014 471134
rect 342545 471218 342781 471454
rect 342545 470898 342781 471134
rect 439581 471218 439817 471454
rect 439581 470898 439817 471134
rect 446517 471218 446753 471454
rect 446517 470898 446753 471134
rect 543553 471218 543789 471454
rect 543553 470898 543789 471134
rect 548058 471218 548294 471454
rect 548378 471218 548614 471454
rect 548058 470898 548294 471134
rect 548378 470898 548614 471134
rect 570292 471218 570528 471454
rect 570612 471218 570848 471454
rect 570292 470898 570528 471134
rect 570612 470898 570848 471134
rect 7876 453218 8112 453454
rect 8196 453218 8432 453454
rect 7876 452898 8112 453134
rect 8196 452898 8432 453134
rect 17658 453218 17894 453454
rect 17978 453218 18214 453454
rect 17658 452898 17894 453134
rect 17978 452898 18214 453134
rect 34897 453218 35133 453454
rect 34897 452898 35133 453134
rect 133373 453218 133609 453454
rect 133373 452898 133609 453134
rect 138869 453218 139105 453454
rect 138869 452898 139105 453134
rect 237345 453218 237581 453454
rect 237345 452898 237581 453134
rect 262458 453218 262694 453454
rect 262778 453218 263014 453454
rect 262458 452898 262694 453134
rect 262778 452898 263014 453134
rect 289658 453218 289894 453454
rect 289978 453218 290214 453454
rect 289658 452898 289894 453134
rect 289978 452898 290214 453134
rect 316858 453218 317094 453454
rect 317178 453218 317414 453454
rect 316858 452898 317094 453134
rect 317178 452898 317414 453134
rect 341825 453218 342061 453454
rect 341825 452898 342061 453134
rect 440301 453218 440537 453454
rect 440301 452898 440537 453134
rect 445797 453218 446033 453454
rect 445797 452898 446033 453134
rect 544273 453218 544509 453454
rect 544273 452898 544509 453134
rect 561658 453218 561894 453454
rect 561978 453218 562214 453454
rect 561658 452898 561894 453134
rect 561978 452898 562214 453134
rect 571532 453218 571768 453454
rect 571852 453218 572088 453454
rect 571532 452898 571768 453134
rect 571852 452898 572088 453134
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect 9116 435218 9352 435454
rect 9436 435218 9672 435454
rect 9116 434898 9352 435134
rect 9436 434898 9672 435134
rect 31258 435218 31494 435454
rect 31578 435218 31814 435454
rect 31258 434898 31494 435134
rect 31578 434898 31814 435134
rect 58458 435218 58694 435454
rect 58778 435218 59014 435454
rect 58458 434898 58694 435134
rect 58778 434898 59014 435134
rect 85658 435218 85894 435454
rect 85978 435218 86214 435454
rect 85658 434898 85894 435134
rect 85978 434898 86214 435134
rect 112858 435218 113094 435454
rect 113178 435218 113414 435454
rect 112858 434898 113094 435134
rect 113178 434898 113414 435134
rect 140058 435218 140294 435454
rect 140378 435218 140614 435454
rect 140058 434898 140294 435134
rect 140378 434898 140614 435134
rect 167258 435218 167494 435454
rect 167578 435218 167814 435454
rect 167258 434898 167494 435134
rect 167578 434898 167814 435134
rect 194458 435218 194694 435454
rect 194778 435218 195014 435454
rect 194458 434898 194694 435134
rect 194778 434898 195014 435134
rect 221658 435218 221894 435454
rect 221978 435218 222214 435454
rect 221658 434898 221894 435134
rect 221978 434898 222214 435134
rect 248858 435218 249094 435454
rect 249178 435218 249414 435454
rect 248858 434898 249094 435134
rect 249178 434898 249414 435134
rect 276058 435218 276294 435454
rect 276378 435218 276614 435454
rect 276058 434898 276294 435134
rect 276378 434898 276614 435134
rect 303258 435218 303494 435454
rect 303578 435218 303814 435454
rect 303258 434898 303494 435134
rect 303578 434898 303814 435134
rect 330458 435218 330694 435454
rect 330778 435218 331014 435454
rect 330458 434898 330694 435134
rect 330778 434898 331014 435134
rect 357658 435218 357894 435454
rect 357978 435218 358214 435454
rect 357658 434898 357894 435134
rect 357978 434898 358214 435134
rect 384858 435218 385094 435454
rect 385178 435218 385414 435454
rect 384858 434898 385094 435134
rect 385178 434898 385414 435134
rect 412058 435218 412294 435454
rect 412378 435218 412614 435454
rect 412058 434898 412294 435134
rect 412378 434898 412614 435134
rect 439258 435218 439494 435454
rect 439578 435218 439814 435454
rect 439258 434898 439494 435134
rect 439578 434898 439814 435134
rect 466458 435218 466694 435454
rect 466778 435218 467014 435454
rect 466458 434898 466694 435134
rect 466778 434898 467014 435134
rect 493658 435218 493894 435454
rect 493978 435218 494214 435454
rect 493658 434898 493894 435134
rect 493978 434898 494214 435134
rect 520858 435218 521094 435454
rect 521178 435218 521414 435454
rect 520858 434898 521094 435134
rect 521178 434898 521414 435134
rect 548058 435218 548294 435454
rect 548378 435218 548614 435454
rect 548058 434898 548294 435134
rect 548378 434898 548614 435134
rect 570292 435218 570528 435454
rect 570612 435218 570848 435454
rect 570292 434898 570528 435134
rect 570612 434898 570848 435134
rect 7876 417218 8112 417454
rect 8196 417218 8432 417454
rect 7876 416898 8112 417134
rect 8196 416898 8432 417134
rect 17658 417218 17894 417454
rect 17978 417218 18214 417454
rect 17658 416898 17894 417134
rect 17978 416898 18214 417134
rect 44858 417218 45094 417454
rect 45178 417218 45414 417454
rect 44858 416898 45094 417134
rect 45178 416898 45414 417134
rect 72058 417218 72294 417454
rect 72378 417218 72614 417454
rect 72058 416898 72294 417134
rect 72378 416898 72614 417134
rect 99258 417218 99494 417454
rect 99578 417218 99814 417454
rect 99258 416898 99494 417134
rect 99578 416898 99814 417134
rect 126458 417218 126694 417454
rect 126778 417218 127014 417454
rect 126458 416898 126694 417134
rect 126778 416898 127014 417134
rect 153658 417218 153894 417454
rect 153978 417218 154214 417454
rect 153658 416898 153894 417134
rect 153978 416898 154214 417134
rect 180858 417218 181094 417454
rect 181178 417218 181414 417454
rect 180858 416898 181094 417134
rect 181178 416898 181414 417134
rect 208058 417218 208294 417454
rect 208378 417218 208614 417454
rect 208058 416898 208294 417134
rect 208378 416898 208614 417134
rect 235258 417218 235494 417454
rect 235578 417218 235814 417454
rect 235258 416898 235494 417134
rect 235578 416898 235814 417134
rect 262458 417218 262694 417454
rect 262778 417218 263014 417454
rect 262458 416898 262694 417134
rect 262778 416898 263014 417134
rect 289658 417218 289894 417454
rect 289978 417218 290214 417454
rect 289658 416898 289894 417134
rect 289978 416898 290214 417134
rect 316858 417218 317094 417454
rect 317178 417218 317414 417454
rect 316858 416898 317094 417134
rect 317178 416898 317414 417134
rect 341825 417218 342061 417454
rect 341825 416898 342061 417134
rect 440301 417218 440537 417454
rect 440301 416898 440537 417134
rect 445797 417218 446033 417454
rect 445797 416898 446033 417134
rect 544273 417218 544509 417454
rect 544273 416898 544509 417134
rect 561658 417218 561894 417454
rect 561978 417218 562214 417454
rect 561658 416898 561894 417134
rect 561978 416898 562214 417134
rect 571532 417218 571768 417454
rect 571852 417218 572088 417454
rect 571532 416898 571768 417134
rect 571852 416898 572088 417134
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect 9116 399218 9352 399454
rect 9436 399218 9672 399454
rect 9116 398898 9352 399134
rect 9436 398898 9672 399134
rect 31258 399218 31494 399454
rect 31578 399218 31814 399454
rect 31258 398898 31494 399134
rect 31578 398898 31814 399134
rect 58458 399218 58694 399454
rect 58778 399218 59014 399454
rect 58458 398898 58694 399134
rect 58778 398898 59014 399134
rect 85658 399218 85894 399454
rect 85978 399218 86214 399454
rect 85658 398898 85894 399134
rect 85978 398898 86214 399134
rect 112858 399218 113094 399454
rect 113178 399218 113414 399454
rect 112858 398898 113094 399134
rect 113178 398898 113414 399134
rect 140058 399218 140294 399454
rect 140378 399218 140614 399454
rect 140058 398898 140294 399134
rect 140378 398898 140614 399134
rect 167258 399218 167494 399454
rect 167578 399218 167814 399454
rect 167258 398898 167494 399134
rect 167578 398898 167814 399134
rect 194458 399218 194694 399454
rect 194778 399218 195014 399454
rect 194458 398898 194694 399134
rect 194778 398898 195014 399134
rect 221658 399218 221894 399454
rect 221978 399218 222214 399454
rect 221658 398898 221894 399134
rect 221978 398898 222214 399134
rect 248858 399218 249094 399454
rect 249178 399218 249414 399454
rect 248858 398898 249094 399134
rect 249178 398898 249414 399134
rect 276058 399218 276294 399454
rect 276378 399218 276614 399454
rect 276058 398898 276294 399134
rect 276378 398898 276614 399134
rect 303258 399218 303494 399454
rect 303578 399218 303814 399454
rect 303258 398898 303494 399134
rect 303578 398898 303814 399134
rect 330458 399218 330694 399454
rect 330778 399218 331014 399454
rect 330458 398898 330694 399134
rect 330778 398898 331014 399134
rect 342545 399218 342781 399454
rect 342545 398898 342781 399134
rect 439581 399218 439817 399454
rect 439581 398898 439817 399134
rect 446517 399218 446753 399454
rect 446517 398898 446753 399134
rect 543553 399218 543789 399454
rect 543553 398898 543789 399134
rect 548058 399218 548294 399454
rect 548378 399218 548614 399454
rect 548058 398898 548294 399134
rect 548378 398898 548614 399134
rect 570292 399218 570528 399454
rect 570612 399218 570848 399454
rect 570292 398898 570528 399134
rect 570612 398898 570848 399134
rect 7876 381218 8112 381454
rect 8196 381218 8432 381454
rect 7876 380898 8112 381134
rect 8196 380898 8432 381134
rect 17658 381218 17894 381454
rect 17978 381218 18214 381454
rect 17658 380898 17894 381134
rect 17978 380898 18214 381134
rect 44858 381218 45094 381454
rect 45178 381218 45414 381454
rect 44858 380898 45094 381134
rect 45178 380898 45414 381134
rect 72058 381218 72294 381454
rect 72378 381218 72614 381454
rect 72058 380898 72294 381134
rect 72378 380898 72614 381134
rect 99258 381218 99494 381454
rect 99578 381218 99814 381454
rect 99258 380898 99494 381134
rect 99578 380898 99814 381134
rect 126458 381218 126694 381454
rect 126778 381218 127014 381454
rect 126458 380898 126694 381134
rect 126778 380898 127014 381134
rect 153658 381218 153894 381454
rect 153978 381218 154214 381454
rect 153658 380898 153894 381134
rect 153978 380898 154214 381134
rect 180858 381218 181094 381454
rect 181178 381218 181414 381454
rect 180858 380898 181094 381134
rect 181178 380898 181414 381134
rect 208058 381218 208294 381454
rect 208378 381218 208614 381454
rect 208058 380898 208294 381134
rect 208378 380898 208614 381134
rect 235258 381218 235494 381454
rect 235578 381218 235814 381454
rect 235258 380898 235494 381134
rect 235578 380898 235814 381134
rect 262458 381218 262694 381454
rect 262778 381218 263014 381454
rect 262458 380898 262694 381134
rect 262778 380898 263014 381134
rect 289658 381218 289894 381454
rect 289978 381218 290214 381454
rect 289658 380898 289894 381134
rect 289978 380898 290214 381134
rect 316858 381218 317094 381454
rect 317178 381218 317414 381454
rect 316858 380898 317094 381134
rect 317178 380898 317414 381134
rect 341825 381218 342061 381454
rect 341825 380898 342061 381134
rect 440301 381218 440537 381454
rect 440301 380898 440537 381134
rect 445797 381218 446033 381454
rect 445797 380898 446033 381134
rect 544273 381218 544509 381454
rect 544273 380898 544509 381134
rect 561658 381218 561894 381454
rect 561978 381218 562214 381454
rect 561658 380898 561894 381134
rect 561978 380898 562214 381134
rect 571532 381218 571768 381454
rect 571852 381218 572088 381454
rect 571532 380898 571768 381134
rect 571852 380898 572088 381134
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect 9116 363218 9352 363454
rect 9436 363218 9672 363454
rect 9116 362898 9352 363134
rect 9436 362898 9672 363134
rect 31258 363218 31494 363454
rect 31578 363218 31814 363454
rect 31258 362898 31494 363134
rect 31578 362898 31814 363134
rect 35617 363218 35853 363454
rect 35617 362898 35853 363134
rect 132653 363218 132889 363454
rect 132653 362898 132889 363134
rect 139589 363218 139825 363454
rect 139589 362898 139825 363134
rect 236625 363218 236861 363454
rect 236625 362898 236861 363134
rect 248858 363218 249094 363454
rect 249178 363218 249414 363454
rect 248858 362898 249094 363134
rect 249178 362898 249414 363134
rect 276058 363218 276294 363454
rect 276378 363218 276614 363454
rect 276058 362898 276294 363134
rect 276378 362898 276614 363134
rect 303258 363218 303494 363454
rect 303578 363218 303814 363454
rect 303258 362898 303494 363134
rect 303578 362898 303814 363134
rect 330458 363218 330694 363454
rect 330778 363218 331014 363454
rect 330458 362898 330694 363134
rect 330778 362898 331014 363134
rect 342545 363218 342781 363454
rect 342545 362898 342781 363134
rect 439581 363218 439817 363454
rect 439581 362898 439817 363134
rect 446517 363218 446753 363454
rect 446517 362898 446753 363134
rect 543553 363218 543789 363454
rect 543553 362898 543789 363134
rect 548058 363218 548294 363454
rect 548378 363218 548614 363454
rect 548058 362898 548294 363134
rect 548378 362898 548614 363134
rect 570292 363218 570528 363454
rect 570612 363218 570848 363454
rect 570292 362898 570528 363134
rect 570612 362898 570848 363134
rect 7876 345218 8112 345454
rect 8196 345218 8432 345454
rect 7876 344898 8112 345134
rect 8196 344898 8432 345134
rect 17658 345218 17894 345454
rect 17978 345218 18214 345454
rect 17658 344898 17894 345134
rect 17978 344898 18214 345134
rect 34897 345218 35133 345454
rect 34897 344898 35133 345134
rect 133373 345218 133609 345454
rect 133373 344898 133609 345134
rect 138869 345218 139105 345454
rect 138869 344898 139105 345134
rect 237345 345218 237581 345454
rect 237345 344898 237581 345134
rect 262458 345218 262694 345454
rect 262778 345218 263014 345454
rect 262458 344898 262694 345134
rect 262778 344898 263014 345134
rect 289658 345218 289894 345454
rect 289978 345218 290214 345454
rect 289658 344898 289894 345134
rect 289978 344898 290214 345134
rect 316858 345218 317094 345454
rect 317178 345218 317414 345454
rect 316858 344898 317094 345134
rect 317178 344898 317414 345134
rect 341825 345218 342061 345454
rect 341825 344898 342061 345134
rect 440301 345218 440537 345454
rect 440301 344898 440537 345134
rect 445797 345218 446033 345454
rect 445797 344898 446033 345134
rect 544273 345218 544509 345454
rect 544273 344898 544509 345134
rect 561658 345218 561894 345454
rect 561978 345218 562214 345454
rect 561658 344898 561894 345134
rect 561978 344898 562214 345134
rect 571532 345218 571768 345454
rect 571852 345218 572088 345454
rect 571532 344898 571768 345134
rect 571852 344898 572088 345134
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect 9116 327218 9352 327454
rect 9436 327218 9672 327454
rect 9116 326898 9352 327134
rect 9436 326898 9672 327134
rect 31258 327218 31494 327454
rect 31578 327218 31814 327454
rect 31258 326898 31494 327134
rect 31578 326898 31814 327134
rect 35617 327218 35853 327454
rect 35617 326898 35853 327134
rect 132653 327218 132889 327454
rect 132653 326898 132889 327134
rect 139589 327218 139825 327454
rect 139589 326898 139825 327134
rect 236625 327218 236861 327454
rect 236625 326898 236861 327134
rect 248858 327218 249094 327454
rect 249178 327218 249414 327454
rect 248858 326898 249094 327134
rect 249178 326898 249414 327134
rect 276058 327218 276294 327454
rect 276378 327218 276614 327454
rect 276058 326898 276294 327134
rect 276378 326898 276614 327134
rect 303258 327218 303494 327454
rect 303578 327218 303814 327454
rect 303258 326898 303494 327134
rect 303578 326898 303814 327134
rect 330458 327218 330694 327454
rect 330778 327218 331014 327454
rect 330458 326898 330694 327134
rect 330778 326898 331014 327134
rect 342545 327218 342781 327454
rect 342545 326898 342781 327134
rect 446517 327218 446753 327454
rect 446517 326898 446753 327134
rect 543553 327218 543789 327454
rect 543553 326898 543789 327134
rect 548058 327218 548294 327454
rect 548378 327218 548614 327454
rect 548058 326898 548294 327134
rect 548378 326898 548614 327134
rect 570292 327218 570528 327454
rect 570612 327218 570848 327454
rect 570292 326898 570528 327134
rect 570612 326898 570848 327134
rect 7876 309218 8112 309454
rect 8196 309218 8432 309454
rect 7876 308898 8112 309134
rect 8196 308898 8432 309134
rect 17658 309218 17894 309454
rect 17978 309218 18214 309454
rect 17658 308898 17894 309134
rect 17978 308898 18214 309134
rect 34897 309218 35133 309454
rect 34897 308898 35133 309134
rect 133373 309218 133609 309454
rect 133373 308898 133609 309134
rect 138869 309218 139105 309454
rect 138869 308898 139105 309134
rect 237345 309218 237581 309454
rect 237345 308898 237581 309134
rect 262458 309218 262694 309454
rect 262778 309218 263014 309454
rect 262458 308898 262694 309134
rect 262778 308898 263014 309134
rect 289658 309218 289894 309454
rect 289978 309218 290214 309454
rect 289658 308898 289894 309134
rect 289978 308898 290214 309134
rect 316858 309218 317094 309454
rect 317178 309218 317414 309454
rect 316858 308898 317094 309134
rect 317178 308898 317414 309134
rect 341825 309218 342061 309454
rect 341825 308898 342061 309134
rect 440301 309218 440537 309454
rect 440301 308898 440537 309134
rect 445797 309218 446033 309454
rect 445797 308898 446033 309134
rect 544273 309218 544509 309454
rect 544273 308898 544509 309134
rect 561658 309218 561894 309454
rect 561978 309218 562214 309454
rect 561658 308898 561894 309134
rect 561978 308898 562214 309134
rect 571532 309218 571768 309454
rect 571852 309218 572088 309454
rect 571532 308898 571768 309134
rect 571852 308898 572088 309134
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect 9116 291218 9352 291454
rect 9436 291218 9672 291454
rect 9116 290898 9352 291134
rect 9436 290898 9672 291134
rect 31258 291218 31494 291454
rect 31578 291218 31814 291454
rect 31258 290898 31494 291134
rect 31578 290898 31814 291134
rect 35617 291218 35853 291454
rect 35617 290898 35853 291134
rect 132653 291218 132889 291454
rect 132653 290898 132889 291134
rect 139589 291218 139825 291454
rect 139589 290898 139825 291134
rect 236625 291218 236861 291454
rect 236625 290898 236861 291134
rect 248858 291218 249094 291454
rect 249178 291218 249414 291454
rect 248858 290898 249094 291134
rect 249178 290898 249414 291134
rect 276058 291218 276294 291454
rect 276378 291218 276614 291454
rect 276058 290898 276294 291134
rect 276378 290898 276614 291134
rect 303258 291218 303494 291454
rect 303578 291218 303814 291454
rect 303258 290898 303494 291134
rect 303578 290898 303814 291134
rect 330458 291218 330694 291454
rect 330778 291218 331014 291454
rect 330458 290898 330694 291134
rect 330778 290898 331014 291134
rect 342545 291218 342781 291454
rect 342545 290898 342781 291134
rect 439581 291218 439817 291454
rect 439581 290898 439817 291134
rect 446517 291218 446753 291454
rect 446517 290898 446753 291134
rect 543553 291218 543789 291454
rect 543553 290898 543789 291134
rect 548058 291218 548294 291454
rect 548378 291218 548614 291454
rect 548058 290898 548294 291134
rect 548378 290898 548614 291134
rect 570292 291218 570528 291454
rect 570612 291218 570848 291454
rect 570292 290898 570528 291134
rect 570612 290898 570848 291134
rect 7876 273218 8112 273454
rect 8196 273218 8432 273454
rect 7876 272898 8112 273134
rect 8196 272898 8432 273134
rect 17658 273218 17894 273454
rect 17978 273218 18214 273454
rect 17658 272898 17894 273134
rect 17978 272898 18214 273134
rect 44858 273218 45094 273454
rect 45178 273218 45414 273454
rect 44858 272898 45094 273134
rect 45178 272898 45414 273134
rect 72058 273218 72294 273454
rect 72378 273218 72614 273454
rect 72058 272898 72294 273134
rect 72378 272898 72614 273134
rect 99258 273218 99494 273454
rect 99578 273218 99814 273454
rect 99258 272898 99494 273134
rect 99578 272898 99814 273134
rect 126458 273218 126694 273454
rect 126778 273218 127014 273454
rect 126458 272898 126694 273134
rect 126778 272898 127014 273134
rect 153658 273218 153894 273454
rect 153978 273218 154214 273454
rect 153658 272898 153894 273134
rect 153978 272898 154214 273134
rect 180858 273218 181094 273454
rect 181178 273218 181414 273454
rect 180858 272898 181094 273134
rect 181178 272898 181414 273134
rect 208058 273218 208294 273454
rect 208378 273218 208614 273454
rect 208058 272898 208294 273134
rect 208378 272898 208614 273134
rect 235258 273218 235494 273454
rect 235578 273218 235814 273454
rect 235258 272898 235494 273134
rect 235578 272898 235814 273134
rect 262458 273218 262694 273454
rect 262778 273218 263014 273454
rect 262458 272898 262694 273134
rect 262778 272898 263014 273134
rect 289658 273218 289894 273454
rect 289978 273218 290214 273454
rect 289658 272898 289894 273134
rect 289978 272898 290214 273134
rect 316858 273218 317094 273454
rect 317178 273218 317414 273454
rect 316858 272898 317094 273134
rect 317178 272898 317414 273134
rect 341825 273218 342061 273454
rect 341825 272898 342061 273134
rect 440301 273218 440537 273454
rect 440301 272898 440537 273134
rect 445797 273218 446033 273454
rect 445797 272898 446033 273134
rect 544273 273218 544509 273454
rect 544273 272898 544509 273134
rect 561658 273218 561894 273454
rect 561978 273218 562214 273454
rect 561658 272898 561894 273134
rect 561978 272898 562214 273134
rect 571532 273218 571768 273454
rect 571852 273218 572088 273454
rect 571532 272898 571768 273134
rect 571852 272898 572088 273134
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect 9116 255218 9352 255454
rect 9436 255218 9672 255454
rect 9116 254898 9352 255134
rect 9436 254898 9672 255134
rect 31258 255218 31494 255454
rect 31578 255218 31814 255454
rect 31258 254898 31494 255134
rect 31578 254898 31814 255134
rect 58458 255218 58694 255454
rect 58778 255218 59014 255454
rect 58458 254898 58694 255134
rect 58778 254898 59014 255134
rect 85658 255218 85894 255454
rect 85978 255218 86214 255454
rect 85658 254898 85894 255134
rect 85978 254898 86214 255134
rect 112858 255218 113094 255454
rect 113178 255218 113414 255454
rect 112858 254898 113094 255134
rect 113178 254898 113414 255134
rect 140058 255218 140294 255454
rect 140378 255218 140614 255454
rect 140058 254898 140294 255134
rect 140378 254898 140614 255134
rect 167258 255218 167494 255454
rect 167578 255218 167814 255454
rect 167258 254898 167494 255134
rect 167578 254898 167814 255134
rect 194458 255218 194694 255454
rect 194778 255218 195014 255454
rect 194458 254898 194694 255134
rect 194778 254898 195014 255134
rect 221658 255218 221894 255454
rect 221978 255218 222214 255454
rect 221658 254898 221894 255134
rect 221978 254898 222214 255134
rect 248858 255218 249094 255454
rect 249178 255218 249414 255454
rect 248858 254898 249094 255134
rect 249178 254898 249414 255134
rect 276058 255218 276294 255454
rect 276378 255218 276614 255454
rect 276058 254898 276294 255134
rect 276378 254898 276614 255134
rect 303258 255218 303494 255454
rect 303578 255218 303814 255454
rect 303258 254898 303494 255134
rect 303578 254898 303814 255134
rect 330458 255218 330694 255454
rect 330778 255218 331014 255454
rect 330458 254898 330694 255134
rect 330778 254898 331014 255134
rect 342545 255218 342781 255454
rect 342545 254898 342781 255134
rect 439581 255218 439817 255454
rect 439581 254898 439817 255134
rect 446517 255218 446753 255454
rect 446517 254898 446753 255134
rect 543553 255218 543789 255454
rect 543553 254898 543789 255134
rect 548058 255218 548294 255454
rect 548378 255218 548614 255454
rect 548058 254898 548294 255134
rect 548378 254898 548614 255134
rect 570292 255218 570528 255454
rect 570612 255218 570848 255454
rect 570292 254898 570528 255134
rect 570612 254898 570848 255134
rect 7876 237218 8112 237454
rect 8196 237218 8432 237454
rect 7876 236898 8112 237134
rect 8196 236898 8432 237134
rect 17658 237218 17894 237454
rect 17978 237218 18214 237454
rect 17658 236898 17894 237134
rect 17978 236898 18214 237134
rect 44858 237218 45094 237454
rect 45178 237218 45414 237454
rect 44858 236898 45094 237134
rect 45178 236898 45414 237134
rect 72058 237218 72294 237454
rect 72378 237218 72614 237454
rect 72058 236898 72294 237134
rect 72378 236898 72614 237134
rect 99258 237218 99494 237454
rect 99578 237218 99814 237454
rect 99258 236898 99494 237134
rect 99578 236898 99814 237134
rect 126458 237218 126694 237454
rect 126778 237218 127014 237454
rect 126458 236898 126694 237134
rect 126778 236898 127014 237134
rect 153658 237218 153894 237454
rect 153978 237218 154214 237454
rect 153658 236898 153894 237134
rect 153978 236898 154214 237134
rect 180858 237218 181094 237454
rect 181178 237218 181414 237454
rect 180858 236898 181094 237134
rect 181178 236898 181414 237134
rect 208058 237218 208294 237454
rect 208378 237218 208614 237454
rect 208058 236898 208294 237134
rect 208378 236898 208614 237134
rect 235258 237218 235494 237454
rect 235578 237218 235814 237454
rect 235258 236898 235494 237134
rect 235578 236898 235814 237134
rect 262458 237218 262694 237454
rect 262778 237218 263014 237454
rect 262458 236898 262694 237134
rect 262778 236898 263014 237134
rect 289658 237218 289894 237454
rect 289978 237218 290214 237454
rect 289658 236898 289894 237134
rect 289978 236898 290214 237134
rect 316858 237218 317094 237454
rect 317178 237218 317414 237454
rect 316858 236898 317094 237134
rect 317178 236898 317414 237134
rect 344058 237218 344294 237454
rect 344378 237218 344614 237454
rect 344058 236898 344294 237134
rect 344378 236898 344614 237134
rect 371258 237218 371494 237454
rect 371578 237218 371814 237454
rect 371258 236898 371494 237134
rect 371578 236898 371814 237134
rect 398458 237218 398694 237454
rect 398778 237218 399014 237454
rect 398458 236898 398694 237134
rect 398778 236898 399014 237134
rect 425658 237218 425894 237454
rect 425978 237218 426214 237454
rect 425658 236898 425894 237134
rect 425978 236898 426214 237134
rect 452858 237218 453094 237454
rect 453178 237218 453414 237454
rect 452858 236898 453094 237134
rect 453178 236898 453414 237134
rect 480058 237218 480294 237454
rect 480378 237218 480614 237454
rect 480058 236898 480294 237134
rect 480378 236898 480614 237134
rect 507258 237218 507494 237454
rect 507578 237218 507814 237454
rect 507258 236898 507494 237134
rect 507578 236898 507814 237134
rect 534458 237218 534694 237454
rect 534778 237218 535014 237454
rect 534458 236898 534694 237134
rect 534778 236898 535014 237134
rect 561658 237218 561894 237454
rect 561978 237218 562214 237454
rect 561658 236898 561894 237134
rect 561978 236898 562214 237134
rect 571532 237218 571768 237454
rect 571852 237218 572088 237454
rect 571532 236898 571768 237134
rect 571852 236898 572088 237134
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect 9116 219218 9352 219454
rect 9436 219218 9672 219454
rect 9116 218898 9352 219134
rect 9436 218898 9672 219134
rect 31258 219218 31494 219454
rect 31578 219218 31814 219454
rect 31258 218898 31494 219134
rect 31578 218898 31814 219134
rect 35617 219218 35853 219454
rect 35617 218898 35853 219134
rect 132653 219218 132889 219454
rect 132653 218898 132889 219134
rect 139589 219218 139825 219454
rect 139589 218898 139825 219134
rect 236625 219218 236861 219454
rect 236625 218898 236861 219134
rect 248858 219218 249094 219454
rect 249178 219218 249414 219454
rect 248858 218898 249094 219134
rect 249178 218898 249414 219134
rect 276058 219218 276294 219454
rect 276378 219218 276614 219454
rect 276058 218898 276294 219134
rect 276378 218898 276614 219134
rect 303258 219218 303494 219454
rect 303578 219218 303814 219454
rect 303258 218898 303494 219134
rect 303578 218898 303814 219134
rect 330458 219218 330694 219454
rect 330778 219218 331014 219454
rect 330458 218898 330694 219134
rect 330778 218898 331014 219134
rect 342545 219218 342781 219454
rect 342545 218898 342781 219134
rect 439581 219218 439817 219454
rect 439581 218898 439817 219134
rect 446517 219218 446753 219454
rect 446517 218898 446753 219134
rect 543553 219218 543789 219454
rect 543553 218898 543789 219134
rect 548058 219218 548294 219454
rect 548378 219218 548614 219454
rect 548058 218898 548294 219134
rect 548378 218898 548614 219134
rect 570292 219218 570528 219454
rect 570612 219218 570848 219454
rect 570292 218898 570528 219134
rect 570612 218898 570848 219134
rect 7876 201218 8112 201454
rect 8196 201218 8432 201454
rect 7876 200898 8112 201134
rect 8196 200898 8432 201134
rect 17658 201218 17894 201454
rect 17978 201218 18214 201454
rect 17658 200898 17894 201134
rect 17978 200898 18214 201134
rect 34897 201218 35133 201454
rect 34897 200898 35133 201134
rect 133373 201218 133609 201454
rect 133373 200898 133609 201134
rect 138869 201218 139105 201454
rect 138869 200898 139105 201134
rect 237345 201218 237581 201454
rect 237345 200898 237581 201134
rect 262458 201218 262694 201454
rect 262778 201218 263014 201454
rect 262458 200898 262694 201134
rect 262778 200898 263014 201134
rect 289658 201218 289894 201454
rect 289978 201218 290214 201454
rect 289658 200898 289894 201134
rect 289978 200898 290214 201134
rect 316858 201218 317094 201454
rect 317178 201218 317414 201454
rect 316858 200898 317094 201134
rect 317178 200898 317414 201134
rect 341825 201218 342061 201454
rect 341825 200898 342061 201134
rect 440301 201218 440537 201454
rect 440301 200898 440537 201134
rect 445797 201218 446033 201454
rect 445797 200898 446033 201134
rect 544273 201218 544509 201454
rect 544273 200898 544509 201134
rect 561658 201218 561894 201454
rect 561978 201218 562214 201454
rect 561658 200898 561894 201134
rect 561978 200898 562214 201134
rect 571532 201218 571768 201454
rect 571852 201218 572088 201454
rect 571532 200898 571768 201134
rect 571852 200898 572088 201134
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect 9116 183218 9352 183454
rect 9436 183218 9672 183454
rect 9116 182898 9352 183134
rect 9436 182898 9672 183134
rect 31258 183218 31494 183454
rect 31578 183218 31814 183454
rect 31258 182898 31494 183134
rect 31578 182898 31814 183134
rect 35617 183218 35853 183454
rect 35617 182898 35853 183134
rect 132653 183218 132889 183454
rect 132653 182898 132889 183134
rect 139589 183218 139825 183454
rect 139589 182898 139825 183134
rect 236625 183218 236861 183454
rect 236625 182898 236861 183134
rect 248858 183218 249094 183454
rect 249178 183218 249414 183454
rect 248858 182898 249094 183134
rect 249178 182898 249414 183134
rect 276058 183218 276294 183454
rect 276378 183218 276614 183454
rect 276058 182898 276294 183134
rect 276378 182898 276614 183134
rect 303258 183218 303494 183454
rect 303578 183218 303814 183454
rect 303258 182898 303494 183134
rect 303578 182898 303814 183134
rect 330458 183218 330694 183454
rect 330778 183218 331014 183454
rect 330458 182898 330694 183134
rect 330778 182898 331014 183134
rect 342545 183218 342781 183454
rect 342545 182898 342781 183134
rect 439581 183218 439817 183454
rect 439581 182898 439817 183134
rect 446517 183218 446753 183454
rect 446517 182898 446753 183134
rect 543553 183218 543789 183454
rect 543553 182898 543789 183134
rect 548058 183218 548294 183454
rect 548378 183218 548614 183454
rect 548058 182898 548294 183134
rect 548378 182898 548614 183134
rect 570292 183218 570528 183454
rect 570612 183218 570848 183454
rect 570292 182898 570528 183134
rect 570612 182898 570848 183134
rect 7876 165218 8112 165454
rect 8196 165218 8432 165454
rect 7876 164898 8112 165134
rect 8196 164898 8432 165134
rect 17658 165218 17894 165454
rect 17978 165218 18214 165454
rect 17658 164898 17894 165134
rect 17978 164898 18214 165134
rect 34897 165218 35133 165454
rect 34897 164898 35133 165134
rect 133373 165218 133609 165454
rect 133373 164898 133609 165134
rect 138869 165218 139105 165454
rect 138869 164898 139105 165134
rect 237345 165218 237581 165454
rect 237345 164898 237581 165134
rect 262458 165218 262694 165454
rect 262778 165218 263014 165454
rect 262458 164898 262694 165134
rect 262778 164898 263014 165134
rect 289658 165218 289894 165454
rect 289978 165218 290214 165454
rect 289658 164898 289894 165134
rect 289978 164898 290214 165134
rect 316858 165218 317094 165454
rect 317178 165218 317414 165454
rect 316858 164898 317094 165134
rect 317178 164898 317414 165134
rect 341825 165218 342061 165454
rect 341825 164898 342061 165134
rect 440301 165218 440537 165454
rect 440301 164898 440537 165134
rect 445797 165218 446033 165454
rect 445797 164898 446033 165134
rect 544273 165218 544509 165454
rect 544273 164898 544509 165134
rect 561658 165218 561894 165454
rect 561978 165218 562214 165454
rect 561658 164898 561894 165134
rect 561978 164898 562214 165134
rect 571532 165218 571768 165454
rect 571852 165218 572088 165454
rect 571532 164898 571768 165134
rect 571852 164898 572088 165134
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect 9116 147218 9352 147454
rect 9436 147218 9672 147454
rect 9116 146898 9352 147134
rect 9436 146898 9672 147134
rect 31258 147218 31494 147454
rect 31578 147218 31814 147454
rect 31258 146898 31494 147134
rect 31578 146898 31814 147134
rect 58458 147218 58694 147454
rect 58778 147218 59014 147454
rect 58458 146898 58694 147134
rect 58778 146898 59014 147134
rect 85658 147218 85894 147454
rect 85978 147218 86214 147454
rect 85658 146898 85894 147134
rect 85978 146898 86214 147134
rect 112858 147218 113094 147454
rect 113178 147218 113414 147454
rect 112858 146898 113094 147134
rect 113178 146898 113414 147134
rect 140058 147218 140294 147454
rect 140378 147218 140614 147454
rect 140058 146898 140294 147134
rect 140378 146898 140614 147134
rect 167258 147218 167494 147454
rect 167578 147218 167814 147454
rect 167258 146898 167494 147134
rect 167578 146898 167814 147134
rect 194458 147218 194694 147454
rect 194778 147218 195014 147454
rect 194458 146898 194694 147134
rect 194778 146898 195014 147134
rect 221658 147218 221894 147454
rect 221978 147218 222214 147454
rect 221658 146898 221894 147134
rect 221978 146898 222214 147134
rect 248858 147218 249094 147454
rect 249178 147218 249414 147454
rect 248858 146898 249094 147134
rect 249178 146898 249414 147134
rect 276058 147218 276294 147454
rect 276378 147218 276614 147454
rect 276058 146898 276294 147134
rect 276378 146898 276614 147134
rect 303258 147218 303494 147454
rect 303578 147218 303814 147454
rect 303258 146898 303494 147134
rect 303578 146898 303814 147134
rect 330458 147218 330694 147454
rect 330778 147218 331014 147454
rect 330458 146898 330694 147134
rect 330778 146898 331014 147134
rect 357658 147218 357894 147454
rect 357978 147218 358214 147454
rect 357658 146898 357894 147134
rect 357978 146898 358214 147134
rect 384858 147218 385094 147454
rect 385178 147218 385414 147454
rect 384858 146898 385094 147134
rect 385178 146898 385414 147134
rect 412058 147218 412294 147454
rect 412378 147218 412614 147454
rect 412058 146898 412294 147134
rect 412378 146898 412614 147134
rect 439258 147218 439494 147454
rect 439578 147218 439814 147454
rect 439258 146898 439494 147134
rect 439578 146898 439814 147134
rect 466458 147218 466694 147454
rect 466778 147218 467014 147454
rect 466458 146898 466694 147134
rect 466778 146898 467014 147134
rect 493658 147218 493894 147454
rect 493978 147218 494214 147454
rect 493658 146898 493894 147134
rect 493978 146898 494214 147134
rect 520858 147218 521094 147454
rect 521178 147218 521414 147454
rect 520858 146898 521094 147134
rect 521178 146898 521414 147134
rect 548058 147218 548294 147454
rect 548378 147218 548614 147454
rect 548058 146898 548294 147134
rect 548378 146898 548614 147134
rect 570292 147218 570528 147454
rect 570612 147218 570848 147454
rect 570292 146898 570528 147134
rect 570612 146898 570848 147134
rect 7876 129218 8112 129454
rect 8196 129218 8432 129454
rect 7876 128898 8112 129134
rect 8196 128898 8432 129134
rect 17658 129218 17894 129454
rect 17978 129218 18214 129454
rect 17658 128898 17894 129134
rect 17978 128898 18214 129134
rect 34897 129218 35133 129454
rect 34897 128898 35133 129134
rect 133373 129218 133609 129454
rect 133373 128898 133609 129134
rect 138869 129218 139105 129454
rect 138869 128898 139105 129134
rect 237345 129218 237581 129454
rect 237345 128898 237581 129134
rect 262458 129218 262694 129454
rect 262778 129218 263014 129454
rect 262458 128898 262694 129134
rect 262778 128898 263014 129134
rect 289658 129218 289894 129454
rect 289978 129218 290214 129454
rect 289658 128898 289894 129134
rect 289978 128898 290214 129134
rect 316858 129218 317094 129454
rect 317178 129218 317414 129454
rect 316858 128898 317094 129134
rect 317178 128898 317414 129134
rect 341825 129218 342061 129454
rect 341825 128898 342061 129134
rect 440301 129218 440537 129454
rect 440301 128898 440537 129134
rect 445797 129218 446033 129454
rect 445797 128898 446033 129134
rect 544273 129218 544509 129454
rect 544273 128898 544509 129134
rect 561658 129218 561894 129454
rect 561978 129218 562214 129454
rect 561658 128898 561894 129134
rect 561978 128898 562214 129134
rect 571532 129218 571768 129454
rect 571852 129218 572088 129454
rect 571532 128898 571768 129134
rect 571852 128898 572088 129134
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect 9116 111218 9352 111454
rect 9436 111218 9672 111454
rect 9116 110898 9352 111134
rect 9436 110898 9672 111134
rect 31258 111218 31494 111454
rect 31578 111218 31814 111454
rect 31258 110898 31494 111134
rect 31578 110898 31814 111134
rect 35617 111218 35853 111454
rect 35617 110898 35853 111134
rect 132653 111218 132889 111454
rect 132653 110898 132889 111134
rect 139589 111218 139825 111454
rect 139589 110898 139825 111134
rect 236625 111218 236861 111454
rect 236625 110898 236861 111134
rect 248858 111218 249094 111454
rect 249178 111218 249414 111454
rect 248858 110898 249094 111134
rect 249178 110898 249414 111134
rect 276058 111218 276294 111454
rect 276378 111218 276614 111454
rect 276058 110898 276294 111134
rect 276378 110898 276614 111134
rect 303258 111218 303494 111454
rect 303578 111218 303814 111454
rect 303258 110898 303494 111134
rect 303578 110898 303814 111134
rect 330458 111218 330694 111454
rect 330778 111218 331014 111454
rect 330458 110898 330694 111134
rect 330778 110898 331014 111134
rect 342545 111218 342781 111454
rect 342545 110898 342781 111134
rect 439581 111218 439817 111454
rect 439581 110898 439817 111134
rect 446517 111218 446753 111454
rect 446517 110898 446753 111134
rect 543553 111218 543789 111454
rect 543553 110898 543789 111134
rect 548058 111218 548294 111454
rect 548378 111218 548614 111454
rect 548058 110898 548294 111134
rect 548378 110898 548614 111134
rect 570292 111218 570528 111454
rect 570612 111218 570848 111454
rect 570292 110898 570528 111134
rect 570612 110898 570848 111134
rect 7876 93218 8112 93454
rect 8196 93218 8432 93454
rect 7876 92898 8112 93134
rect 8196 92898 8432 93134
rect 17658 93218 17894 93454
rect 17978 93218 18214 93454
rect 17658 92898 17894 93134
rect 17978 92898 18214 93134
rect 34897 93218 35133 93454
rect 34897 92898 35133 93134
rect 133373 93218 133609 93454
rect 133373 92898 133609 93134
rect 138869 93218 139105 93454
rect 138869 92898 139105 93134
rect 237345 93218 237581 93454
rect 237345 92898 237581 93134
rect 262458 93218 262694 93454
rect 262778 93218 263014 93454
rect 262458 92898 262694 93134
rect 262778 92898 263014 93134
rect 289658 93218 289894 93454
rect 289978 93218 290214 93454
rect 289658 92898 289894 93134
rect 289978 92898 290214 93134
rect 316858 93218 317094 93454
rect 317178 93218 317414 93454
rect 316858 92898 317094 93134
rect 317178 92898 317414 93134
rect 341825 93218 342061 93454
rect 341825 92898 342061 93134
rect 440301 93218 440537 93454
rect 440301 92898 440537 93134
rect 445797 93218 446033 93454
rect 445797 92898 446033 93134
rect 544273 93218 544509 93454
rect 544273 92898 544509 93134
rect 561658 93218 561894 93454
rect 561978 93218 562214 93454
rect 561658 92898 561894 93134
rect 561978 92898 562214 93134
rect 571532 93218 571768 93454
rect 571852 93218 572088 93454
rect 571532 92898 571768 93134
rect 571852 92898 572088 93134
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect 9116 75218 9352 75454
rect 9436 75218 9672 75454
rect 9116 74898 9352 75134
rect 9436 74898 9672 75134
rect 31258 75218 31494 75454
rect 31578 75218 31814 75454
rect 31258 74898 31494 75134
rect 31578 74898 31814 75134
rect 35617 75218 35853 75454
rect 35617 74898 35853 75134
rect 132653 75218 132889 75454
rect 132653 74898 132889 75134
rect 139589 75218 139825 75454
rect 139589 74898 139825 75134
rect 236625 75218 236861 75454
rect 236625 74898 236861 75134
rect 248858 75218 249094 75454
rect 249178 75218 249414 75454
rect 248858 74898 249094 75134
rect 249178 74898 249414 75134
rect 276058 75218 276294 75454
rect 276378 75218 276614 75454
rect 276058 74898 276294 75134
rect 276378 74898 276614 75134
rect 303258 75218 303494 75454
rect 303578 75218 303814 75454
rect 303258 74898 303494 75134
rect 303578 74898 303814 75134
rect 330458 75218 330694 75454
rect 330778 75218 331014 75454
rect 330458 74898 330694 75134
rect 330778 74898 331014 75134
rect 342545 75218 342781 75454
rect 342545 74898 342781 75134
rect 439581 75218 439817 75454
rect 439581 74898 439817 75134
rect 446517 75218 446753 75454
rect 446517 74898 446753 75134
rect 543553 75218 543789 75454
rect 543553 74898 543789 75134
rect 548058 75218 548294 75454
rect 548378 75218 548614 75454
rect 548058 74898 548294 75134
rect 548378 74898 548614 75134
rect 570292 75218 570528 75454
rect 570612 75218 570848 75454
rect 570292 74898 570528 75134
rect 570612 74898 570848 75134
rect 7876 57218 8112 57454
rect 8196 57218 8432 57454
rect 7876 56898 8112 57134
rect 8196 56898 8432 57134
rect 17658 57218 17894 57454
rect 17978 57218 18214 57454
rect 17658 56898 17894 57134
rect 17978 56898 18214 57134
rect 34897 57218 35133 57454
rect 34897 56898 35133 57134
rect 133373 57218 133609 57454
rect 133373 56898 133609 57134
rect 138869 57218 139105 57454
rect 138869 56898 139105 57134
rect 237345 57218 237581 57454
rect 237345 56898 237581 57134
rect 262458 57218 262694 57454
rect 262778 57218 263014 57454
rect 262458 56898 262694 57134
rect 262778 56898 263014 57134
rect 289658 57218 289894 57454
rect 289978 57218 290214 57454
rect 289658 56898 289894 57134
rect 289978 56898 290214 57134
rect 316858 57218 317094 57454
rect 317178 57218 317414 57454
rect 316858 56898 317094 57134
rect 317178 56898 317414 57134
rect 341825 57218 342061 57454
rect 341825 56898 342061 57134
rect 440301 57218 440537 57454
rect 440301 56898 440537 57134
rect 445797 57218 446033 57454
rect 445797 56898 446033 57134
rect 544273 57218 544509 57454
rect 544273 56898 544509 57134
rect 561658 57218 561894 57454
rect 561978 57218 562214 57454
rect 561658 56898 561894 57134
rect 561978 56898 562214 57134
rect 571532 57218 571768 57454
rect 571852 57218 572088 57454
rect 571532 56898 571768 57134
rect 571852 56898 572088 57134
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect 9116 39218 9352 39454
rect 9436 39218 9672 39454
rect 9116 38898 9352 39134
rect 9436 38898 9672 39134
rect 31258 39218 31494 39454
rect 31578 39218 31814 39454
rect 31258 38898 31494 39134
rect 31578 38898 31814 39134
rect 58458 39218 58694 39454
rect 58778 39218 59014 39454
rect 58458 38898 58694 39134
rect 58778 38898 59014 39134
rect 85658 39218 85894 39454
rect 85978 39218 86214 39454
rect 85658 38898 85894 39134
rect 85978 38898 86214 39134
rect 112858 39218 113094 39454
rect 113178 39218 113414 39454
rect 112858 38898 113094 39134
rect 113178 38898 113414 39134
rect 140058 39218 140294 39454
rect 140378 39218 140614 39454
rect 140058 38898 140294 39134
rect 140378 38898 140614 39134
rect 167258 39218 167494 39454
rect 167578 39218 167814 39454
rect 167258 38898 167494 39134
rect 167578 38898 167814 39134
rect 194458 39218 194694 39454
rect 194778 39218 195014 39454
rect 194458 38898 194694 39134
rect 194778 38898 195014 39134
rect 221658 39218 221894 39454
rect 221978 39218 222214 39454
rect 221658 38898 221894 39134
rect 221978 38898 222214 39134
rect 248858 39218 249094 39454
rect 249178 39218 249414 39454
rect 248858 38898 249094 39134
rect 249178 38898 249414 39134
rect 276058 39218 276294 39454
rect 276378 39218 276614 39454
rect 276058 38898 276294 39134
rect 276378 38898 276614 39134
rect 303258 39218 303494 39454
rect 303578 39218 303814 39454
rect 303258 38898 303494 39134
rect 303578 38898 303814 39134
rect 330458 39218 330694 39454
rect 330778 39218 331014 39454
rect 330458 38898 330694 39134
rect 330778 38898 331014 39134
rect 357658 39218 357894 39454
rect 357978 39218 358214 39454
rect 357658 38898 357894 39134
rect 357978 38898 358214 39134
rect 384858 39218 385094 39454
rect 385178 39218 385414 39454
rect 384858 38898 385094 39134
rect 385178 38898 385414 39134
rect 412058 39218 412294 39454
rect 412378 39218 412614 39454
rect 412058 38898 412294 39134
rect 412378 38898 412614 39134
rect 439258 39218 439494 39454
rect 439578 39218 439814 39454
rect 439258 38898 439494 39134
rect 439578 38898 439814 39134
rect 466458 39218 466694 39454
rect 466778 39218 467014 39454
rect 466458 38898 466694 39134
rect 466778 38898 467014 39134
rect 493658 39218 493894 39454
rect 493978 39218 494214 39454
rect 493658 38898 493894 39134
rect 493978 38898 494214 39134
rect 520858 39218 521094 39454
rect 521178 39218 521414 39454
rect 520858 38898 521094 39134
rect 521178 38898 521414 39134
rect 548058 39218 548294 39454
rect 548378 39218 548614 39454
rect 548058 38898 548294 39134
rect 548378 38898 548614 39134
rect 570292 39218 570528 39454
rect 570612 39218 570848 39454
rect 570292 38898 570528 39134
rect 570612 38898 570848 39134
rect 7876 21218 8112 21454
rect 8196 21218 8432 21454
rect 7876 20898 8112 21134
rect 8196 20898 8432 21134
rect 17658 21218 17894 21454
rect 17978 21218 18214 21454
rect 17658 20898 17894 21134
rect 17978 20898 18214 21134
rect 44858 21218 45094 21454
rect 45178 21218 45414 21454
rect 44858 20898 45094 21134
rect 45178 20898 45414 21134
rect 72058 21218 72294 21454
rect 72378 21218 72614 21454
rect 72058 20898 72294 21134
rect 72378 20898 72614 21134
rect 99258 21218 99494 21454
rect 99578 21218 99814 21454
rect 99258 20898 99494 21134
rect 99578 20898 99814 21134
rect 126458 21218 126694 21454
rect 126778 21218 127014 21454
rect 126458 20898 126694 21134
rect 126778 20898 127014 21134
rect 153658 21218 153894 21454
rect 153978 21218 154214 21454
rect 153658 20898 153894 21134
rect 153978 20898 154214 21134
rect 180858 21218 181094 21454
rect 181178 21218 181414 21454
rect 180858 20898 181094 21134
rect 181178 20898 181414 21134
rect 208058 21218 208294 21454
rect 208378 21218 208614 21454
rect 208058 20898 208294 21134
rect 208378 20898 208614 21134
rect 235258 21218 235494 21454
rect 235578 21218 235814 21454
rect 235258 20898 235494 21134
rect 235578 20898 235814 21134
rect 262458 21218 262694 21454
rect 262778 21218 263014 21454
rect 262458 20898 262694 21134
rect 262778 20898 263014 21134
rect 289658 21218 289894 21454
rect 289978 21218 290214 21454
rect 289658 20898 289894 21134
rect 289978 20898 290214 21134
rect 316858 21218 317094 21454
rect 317178 21218 317414 21454
rect 316858 20898 317094 21134
rect 317178 20898 317414 21134
rect 344058 21218 344294 21454
rect 344378 21218 344614 21454
rect 344058 20898 344294 21134
rect 344378 20898 344614 21134
rect 371258 21218 371494 21454
rect 371578 21218 371814 21454
rect 371258 20898 371494 21134
rect 371578 20898 371814 21134
rect 398458 21218 398694 21454
rect 398778 21218 399014 21454
rect 398458 20898 398694 21134
rect 398778 20898 399014 21134
rect 425658 21218 425894 21454
rect 425978 21218 426214 21454
rect 425658 20898 425894 21134
rect 425978 20898 426214 21134
rect 452858 21218 453094 21454
rect 453178 21218 453414 21454
rect 452858 20898 453094 21134
rect 453178 20898 453414 21134
rect 480058 21218 480294 21454
rect 480378 21218 480614 21454
rect 480058 20898 480294 21134
rect 480378 20898 480614 21134
rect 507258 21218 507494 21454
rect 507578 21218 507814 21454
rect 507258 20898 507494 21134
rect 507578 20898 507814 21134
rect 534458 21218 534694 21454
rect 534778 21218 535014 21454
rect 534458 20898 534694 21134
rect 534778 20898 535014 21134
rect 561658 21218 561894 21454
rect 561978 21218 562214 21454
rect 561658 20898 561894 21134
rect 561978 20898 562214 21134
rect 571532 21218 571768 21454
rect 571852 21218 572088 21454
rect 571532 20898 571768 21134
rect 571852 20898 572088 21134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 9116 687454
rect 9352 687218 9436 687454
rect 9672 687218 31258 687454
rect 31494 687218 31578 687454
rect 31814 687218 58458 687454
rect 58694 687218 58778 687454
rect 59014 687218 85658 687454
rect 85894 687218 85978 687454
rect 86214 687218 112858 687454
rect 113094 687218 113178 687454
rect 113414 687218 140058 687454
rect 140294 687218 140378 687454
rect 140614 687218 167258 687454
rect 167494 687218 167578 687454
rect 167814 687218 194458 687454
rect 194694 687218 194778 687454
rect 195014 687218 221658 687454
rect 221894 687218 221978 687454
rect 222214 687218 248858 687454
rect 249094 687218 249178 687454
rect 249414 687218 276058 687454
rect 276294 687218 276378 687454
rect 276614 687218 303258 687454
rect 303494 687218 303578 687454
rect 303814 687218 330458 687454
rect 330694 687218 330778 687454
rect 331014 687218 357658 687454
rect 357894 687218 357978 687454
rect 358214 687218 384858 687454
rect 385094 687218 385178 687454
rect 385414 687218 412058 687454
rect 412294 687218 412378 687454
rect 412614 687218 439258 687454
rect 439494 687218 439578 687454
rect 439814 687218 466458 687454
rect 466694 687218 466778 687454
rect 467014 687218 493658 687454
rect 493894 687218 493978 687454
rect 494214 687218 520858 687454
rect 521094 687218 521178 687454
rect 521414 687218 548058 687454
rect 548294 687218 548378 687454
rect 548614 687218 570292 687454
rect 570528 687218 570612 687454
rect 570848 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 9116 687134
rect 9352 686898 9436 687134
rect 9672 686898 31258 687134
rect 31494 686898 31578 687134
rect 31814 686898 58458 687134
rect 58694 686898 58778 687134
rect 59014 686898 85658 687134
rect 85894 686898 85978 687134
rect 86214 686898 112858 687134
rect 113094 686898 113178 687134
rect 113414 686898 140058 687134
rect 140294 686898 140378 687134
rect 140614 686898 167258 687134
rect 167494 686898 167578 687134
rect 167814 686898 194458 687134
rect 194694 686898 194778 687134
rect 195014 686898 221658 687134
rect 221894 686898 221978 687134
rect 222214 686898 248858 687134
rect 249094 686898 249178 687134
rect 249414 686898 276058 687134
rect 276294 686898 276378 687134
rect 276614 686898 303258 687134
rect 303494 686898 303578 687134
rect 303814 686898 330458 687134
rect 330694 686898 330778 687134
rect 331014 686898 357658 687134
rect 357894 686898 357978 687134
rect 358214 686898 384858 687134
rect 385094 686898 385178 687134
rect 385414 686898 412058 687134
rect 412294 686898 412378 687134
rect 412614 686898 439258 687134
rect 439494 686898 439578 687134
rect 439814 686898 466458 687134
rect 466694 686898 466778 687134
rect 467014 686898 493658 687134
rect 493894 686898 493978 687134
rect 494214 686898 520858 687134
rect 521094 686898 521178 687134
rect 521414 686898 548058 687134
rect 548294 686898 548378 687134
rect 548614 686898 570292 687134
rect 570528 686898 570612 687134
rect 570848 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 7876 669454
rect 8112 669218 8196 669454
rect 8432 669218 17658 669454
rect 17894 669218 17978 669454
rect 18214 669218 44858 669454
rect 45094 669218 45178 669454
rect 45414 669218 72058 669454
rect 72294 669218 72378 669454
rect 72614 669218 99258 669454
rect 99494 669218 99578 669454
rect 99814 669218 126458 669454
rect 126694 669218 126778 669454
rect 127014 669218 153658 669454
rect 153894 669218 153978 669454
rect 154214 669218 180858 669454
rect 181094 669218 181178 669454
rect 181414 669218 208058 669454
rect 208294 669218 208378 669454
rect 208614 669218 235258 669454
rect 235494 669218 235578 669454
rect 235814 669218 262458 669454
rect 262694 669218 262778 669454
rect 263014 669218 289658 669454
rect 289894 669218 289978 669454
rect 290214 669218 316858 669454
rect 317094 669218 317178 669454
rect 317414 669218 344058 669454
rect 344294 669218 344378 669454
rect 344614 669218 371258 669454
rect 371494 669218 371578 669454
rect 371814 669218 398458 669454
rect 398694 669218 398778 669454
rect 399014 669218 425658 669454
rect 425894 669218 425978 669454
rect 426214 669218 452858 669454
rect 453094 669218 453178 669454
rect 453414 669218 480058 669454
rect 480294 669218 480378 669454
rect 480614 669218 507258 669454
rect 507494 669218 507578 669454
rect 507814 669218 534458 669454
rect 534694 669218 534778 669454
rect 535014 669218 561658 669454
rect 561894 669218 561978 669454
rect 562214 669218 571532 669454
rect 571768 669218 571852 669454
rect 572088 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 7876 669134
rect 8112 668898 8196 669134
rect 8432 668898 17658 669134
rect 17894 668898 17978 669134
rect 18214 668898 44858 669134
rect 45094 668898 45178 669134
rect 45414 668898 72058 669134
rect 72294 668898 72378 669134
rect 72614 668898 99258 669134
rect 99494 668898 99578 669134
rect 99814 668898 126458 669134
rect 126694 668898 126778 669134
rect 127014 668898 153658 669134
rect 153894 668898 153978 669134
rect 154214 668898 180858 669134
rect 181094 668898 181178 669134
rect 181414 668898 208058 669134
rect 208294 668898 208378 669134
rect 208614 668898 235258 669134
rect 235494 668898 235578 669134
rect 235814 668898 262458 669134
rect 262694 668898 262778 669134
rect 263014 668898 289658 669134
rect 289894 668898 289978 669134
rect 290214 668898 316858 669134
rect 317094 668898 317178 669134
rect 317414 668898 344058 669134
rect 344294 668898 344378 669134
rect 344614 668898 371258 669134
rect 371494 668898 371578 669134
rect 371814 668898 398458 669134
rect 398694 668898 398778 669134
rect 399014 668898 425658 669134
rect 425894 668898 425978 669134
rect 426214 668898 452858 669134
rect 453094 668898 453178 669134
rect 453414 668898 480058 669134
rect 480294 668898 480378 669134
rect 480614 668898 507258 669134
rect 507494 668898 507578 669134
rect 507814 668898 534458 669134
rect 534694 668898 534778 669134
rect 535014 668898 561658 669134
rect 561894 668898 561978 669134
rect 562214 668898 571532 669134
rect 571768 668898 571852 669134
rect 572088 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 9116 651454
rect 9352 651218 9436 651454
rect 9672 651218 31258 651454
rect 31494 651218 31578 651454
rect 31814 651218 58458 651454
rect 58694 651218 58778 651454
rect 59014 651218 85658 651454
rect 85894 651218 85978 651454
rect 86214 651218 112858 651454
rect 113094 651218 113178 651454
rect 113414 651218 140058 651454
rect 140294 651218 140378 651454
rect 140614 651218 167258 651454
rect 167494 651218 167578 651454
rect 167814 651218 194458 651454
rect 194694 651218 194778 651454
rect 195014 651218 221658 651454
rect 221894 651218 221978 651454
rect 222214 651218 248858 651454
rect 249094 651218 249178 651454
rect 249414 651218 276058 651454
rect 276294 651218 276378 651454
rect 276614 651218 303258 651454
rect 303494 651218 303578 651454
rect 303814 651218 330458 651454
rect 330694 651218 330778 651454
rect 331014 651218 357658 651454
rect 357894 651218 357978 651454
rect 358214 651218 384858 651454
rect 385094 651218 385178 651454
rect 385414 651218 412058 651454
rect 412294 651218 412378 651454
rect 412614 651218 439258 651454
rect 439494 651218 439578 651454
rect 439814 651218 466458 651454
rect 466694 651218 466778 651454
rect 467014 651218 493658 651454
rect 493894 651218 493978 651454
rect 494214 651218 520858 651454
rect 521094 651218 521178 651454
rect 521414 651218 548058 651454
rect 548294 651218 548378 651454
rect 548614 651218 570292 651454
rect 570528 651218 570612 651454
rect 570848 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 9116 651134
rect 9352 650898 9436 651134
rect 9672 650898 31258 651134
rect 31494 650898 31578 651134
rect 31814 650898 58458 651134
rect 58694 650898 58778 651134
rect 59014 650898 85658 651134
rect 85894 650898 85978 651134
rect 86214 650898 112858 651134
rect 113094 650898 113178 651134
rect 113414 650898 140058 651134
rect 140294 650898 140378 651134
rect 140614 650898 167258 651134
rect 167494 650898 167578 651134
rect 167814 650898 194458 651134
rect 194694 650898 194778 651134
rect 195014 650898 221658 651134
rect 221894 650898 221978 651134
rect 222214 650898 248858 651134
rect 249094 650898 249178 651134
rect 249414 650898 276058 651134
rect 276294 650898 276378 651134
rect 276614 650898 303258 651134
rect 303494 650898 303578 651134
rect 303814 650898 330458 651134
rect 330694 650898 330778 651134
rect 331014 650898 357658 651134
rect 357894 650898 357978 651134
rect 358214 650898 384858 651134
rect 385094 650898 385178 651134
rect 385414 650898 412058 651134
rect 412294 650898 412378 651134
rect 412614 650898 439258 651134
rect 439494 650898 439578 651134
rect 439814 650898 466458 651134
rect 466694 650898 466778 651134
rect 467014 650898 493658 651134
rect 493894 650898 493978 651134
rect 494214 650898 520858 651134
rect 521094 650898 521178 651134
rect 521414 650898 548058 651134
rect 548294 650898 548378 651134
rect 548614 650898 570292 651134
rect 570528 650898 570612 651134
rect 570848 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 7876 633454
rect 8112 633218 8196 633454
rect 8432 633218 17658 633454
rect 17894 633218 17978 633454
rect 18214 633218 44858 633454
rect 45094 633218 45178 633454
rect 45414 633218 72058 633454
rect 72294 633218 72378 633454
rect 72614 633218 99258 633454
rect 99494 633218 99578 633454
rect 99814 633218 126458 633454
rect 126694 633218 126778 633454
rect 127014 633218 153658 633454
rect 153894 633218 153978 633454
rect 154214 633218 180858 633454
rect 181094 633218 181178 633454
rect 181414 633218 208058 633454
rect 208294 633218 208378 633454
rect 208614 633218 235258 633454
rect 235494 633218 235578 633454
rect 235814 633218 262458 633454
rect 262694 633218 262778 633454
rect 263014 633218 289658 633454
rect 289894 633218 289978 633454
rect 290214 633218 316858 633454
rect 317094 633218 317178 633454
rect 317414 633218 344058 633454
rect 344294 633218 344378 633454
rect 344614 633218 371258 633454
rect 371494 633218 371578 633454
rect 371814 633218 398458 633454
rect 398694 633218 398778 633454
rect 399014 633218 425658 633454
rect 425894 633218 425978 633454
rect 426214 633218 452858 633454
rect 453094 633218 453178 633454
rect 453414 633218 480058 633454
rect 480294 633218 480378 633454
rect 480614 633218 507258 633454
rect 507494 633218 507578 633454
rect 507814 633218 534458 633454
rect 534694 633218 534778 633454
rect 535014 633218 561658 633454
rect 561894 633218 561978 633454
rect 562214 633218 571532 633454
rect 571768 633218 571852 633454
rect 572088 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 7876 633134
rect 8112 632898 8196 633134
rect 8432 632898 17658 633134
rect 17894 632898 17978 633134
rect 18214 632898 44858 633134
rect 45094 632898 45178 633134
rect 45414 632898 72058 633134
rect 72294 632898 72378 633134
rect 72614 632898 99258 633134
rect 99494 632898 99578 633134
rect 99814 632898 126458 633134
rect 126694 632898 126778 633134
rect 127014 632898 153658 633134
rect 153894 632898 153978 633134
rect 154214 632898 180858 633134
rect 181094 632898 181178 633134
rect 181414 632898 208058 633134
rect 208294 632898 208378 633134
rect 208614 632898 235258 633134
rect 235494 632898 235578 633134
rect 235814 632898 262458 633134
rect 262694 632898 262778 633134
rect 263014 632898 289658 633134
rect 289894 632898 289978 633134
rect 290214 632898 316858 633134
rect 317094 632898 317178 633134
rect 317414 632898 344058 633134
rect 344294 632898 344378 633134
rect 344614 632898 371258 633134
rect 371494 632898 371578 633134
rect 371814 632898 398458 633134
rect 398694 632898 398778 633134
rect 399014 632898 425658 633134
rect 425894 632898 425978 633134
rect 426214 632898 452858 633134
rect 453094 632898 453178 633134
rect 453414 632898 480058 633134
rect 480294 632898 480378 633134
rect 480614 632898 507258 633134
rect 507494 632898 507578 633134
rect 507814 632898 534458 633134
rect 534694 632898 534778 633134
rect 535014 632898 561658 633134
rect 561894 632898 561978 633134
rect 562214 632898 571532 633134
rect 571768 632898 571852 633134
rect 572088 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 9116 615454
rect 9352 615218 9436 615454
rect 9672 615218 31258 615454
rect 31494 615218 31578 615454
rect 31814 615218 58458 615454
rect 58694 615218 58778 615454
rect 59014 615218 85658 615454
rect 85894 615218 85978 615454
rect 86214 615218 112858 615454
rect 113094 615218 113178 615454
rect 113414 615218 140058 615454
rect 140294 615218 140378 615454
rect 140614 615218 167258 615454
rect 167494 615218 167578 615454
rect 167814 615218 194458 615454
rect 194694 615218 194778 615454
rect 195014 615218 221658 615454
rect 221894 615218 221978 615454
rect 222214 615218 248858 615454
rect 249094 615218 249178 615454
rect 249414 615218 276058 615454
rect 276294 615218 276378 615454
rect 276614 615218 303258 615454
rect 303494 615218 303578 615454
rect 303814 615218 330458 615454
rect 330694 615218 330778 615454
rect 331014 615218 357658 615454
rect 357894 615218 357978 615454
rect 358214 615218 384858 615454
rect 385094 615218 385178 615454
rect 385414 615218 412058 615454
rect 412294 615218 412378 615454
rect 412614 615218 439258 615454
rect 439494 615218 439578 615454
rect 439814 615218 466458 615454
rect 466694 615218 466778 615454
rect 467014 615218 493658 615454
rect 493894 615218 493978 615454
rect 494214 615218 520858 615454
rect 521094 615218 521178 615454
rect 521414 615218 548058 615454
rect 548294 615218 548378 615454
rect 548614 615218 570292 615454
rect 570528 615218 570612 615454
rect 570848 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 9116 615134
rect 9352 614898 9436 615134
rect 9672 614898 31258 615134
rect 31494 614898 31578 615134
rect 31814 614898 58458 615134
rect 58694 614898 58778 615134
rect 59014 614898 85658 615134
rect 85894 614898 85978 615134
rect 86214 614898 112858 615134
rect 113094 614898 113178 615134
rect 113414 614898 140058 615134
rect 140294 614898 140378 615134
rect 140614 614898 167258 615134
rect 167494 614898 167578 615134
rect 167814 614898 194458 615134
rect 194694 614898 194778 615134
rect 195014 614898 221658 615134
rect 221894 614898 221978 615134
rect 222214 614898 248858 615134
rect 249094 614898 249178 615134
rect 249414 614898 276058 615134
rect 276294 614898 276378 615134
rect 276614 614898 303258 615134
rect 303494 614898 303578 615134
rect 303814 614898 330458 615134
rect 330694 614898 330778 615134
rect 331014 614898 357658 615134
rect 357894 614898 357978 615134
rect 358214 614898 384858 615134
rect 385094 614898 385178 615134
rect 385414 614898 412058 615134
rect 412294 614898 412378 615134
rect 412614 614898 439258 615134
rect 439494 614898 439578 615134
rect 439814 614898 466458 615134
rect 466694 614898 466778 615134
rect 467014 614898 493658 615134
rect 493894 614898 493978 615134
rect 494214 614898 520858 615134
rect 521094 614898 521178 615134
rect 521414 614898 548058 615134
rect 548294 614898 548378 615134
rect 548614 614898 570292 615134
rect 570528 614898 570612 615134
rect 570848 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 7876 597454
rect 8112 597218 8196 597454
rect 8432 597218 17658 597454
rect 17894 597218 17978 597454
rect 18214 597218 34897 597454
rect 35133 597218 133373 597454
rect 133609 597218 138869 597454
rect 139105 597218 237345 597454
rect 237581 597218 262458 597454
rect 262694 597218 262778 597454
rect 263014 597218 289658 597454
rect 289894 597218 289978 597454
rect 290214 597218 316858 597454
rect 317094 597218 317178 597454
rect 317414 597218 341825 597454
rect 342061 597218 440301 597454
rect 440537 597218 445797 597454
rect 446033 597218 544273 597454
rect 544509 597218 561658 597454
rect 561894 597218 561978 597454
rect 562214 597218 571532 597454
rect 571768 597218 571852 597454
rect 572088 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 7876 597134
rect 8112 596898 8196 597134
rect 8432 596898 17658 597134
rect 17894 596898 17978 597134
rect 18214 596898 34897 597134
rect 35133 596898 133373 597134
rect 133609 596898 138869 597134
rect 139105 596898 237345 597134
rect 237581 596898 262458 597134
rect 262694 596898 262778 597134
rect 263014 596898 289658 597134
rect 289894 596898 289978 597134
rect 290214 596898 316858 597134
rect 317094 596898 317178 597134
rect 317414 596898 341825 597134
rect 342061 596898 440301 597134
rect 440537 596898 445797 597134
rect 446033 596898 544273 597134
rect 544509 596898 561658 597134
rect 561894 596898 561978 597134
rect 562214 596898 571532 597134
rect 571768 596898 571852 597134
rect 572088 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 9116 579454
rect 9352 579218 9436 579454
rect 9672 579218 31258 579454
rect 31494 579218 31578 579454
rect 31814 579218 35617 579454
rect 35853 579218 132653 579454
rect 132889 579218 139589 579454
rect 139825 579218 236625 579454
rect 236861 579218 248858 579454
rect 249094 579218 249178 579454
rect 249414 579218 276058 579454
rect 276294 579218 276378 579454
rect 276614 579218 303258 579454
rect 303494 579218 303578 579454
rect 303814 579218 330458 579454
rect 330694 579218 330778 579454
rect 331014 579218 342545 579454
rect 342781 579218 439581 579454
rect 439817 579218 446517 579454
rect 446753 579218 543553 579454
rect 543789 579218 548058 579454
rect 548294 579218 548378 579454
rect 548614 579218 570292 579454
rect 570528 579218 570612 579454
rect 570848 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 9116 579134
rect 9352 578898 9436 579134
rect 9672 578898 31258 579134
rect 31494 578898 31578 579134
rect 31814 578898 35617 579134
rect 35853 578898 132653 579134
rect 132889 578898 139589 579134
rect 139825 578898 236625 579134
rect 236861 578898 248858 579134
rect 249094 578898 249178 579134
rect 249414 578898 276058 579134
rect 276294 578898 276378 579134
rect 276614 578898 303258 579134
rect 303494 578898 303578 579134
rect 303814 578898 330458 579134
rect 330694 578898 330778 579134
rect 331014 578898 342545 579134
rect 342781 578898 439581 579134
rect 439817 578898 446517 579134
rect 446753 578898 543553 579134
rect 543789 578898 548058 579134
rect 548294 578898 548378 579134
rect 548614 578898 570292 579134
rect 570528 578898 570612 579134
rect 570848 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 7876 561454
rect 8112 561218 8196 561454
rect 8432 561218 17658 561454
rect 17894 561218 17978 561454
rect 18214 561218 34897 561454
rect 35133 561218 133373 561454
rect 133609 561218 138869 561454
rect 139105 561218 237345 561454
rect 237581 561218 262458 561454
rect 262694 561218 262778 561454
rect 263014 561218 289658 561454
rect 289894 561218 289978 561454
rect 290214 561218 316858 561454
rect 317094 561218 317178 561454
rect 317414 561218 341825 561454
rect 342061 561218 440301 561454
rect 440537 561218 445797 561454
rect 446033 561218 544273 561454
rect 544509 561218 561658 561454
rect 561894 561218 561978 561454
rect 562214 561218 571532 561454
rect 571768 561218 571852 561454
rect 572088 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 7876 561134
rect 8112 560898 8196 561134
rect 8432 560898 17658 561134
rect 17894 560898 17978 561134
rect 18214 560898 34897 561134
rect 35133 560898 133373 561134
rect 133609 560898 138869 561134
rect 139105 560898 237345 561134
rect 237581 560898 262458 561134
rect 262694 560898 262778 561134
rect 263014 560898 289658 561134
rect 289894 560898 289978 561134
rect 290214 560898 316858 561134
rect 317094 560898 317178 561134
rect 317414 560898 341825 561134
rect 342061 560898 440301 561134
rect 440537 560898 445797 561134
rect 446033 560898 544273 561134
rect 544509 560898 561658 561134
rect 561894 560898 561978 561134
rect 562214 560898 571532 561134
rect 571768 560898 571852 561134
rect 572088 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 9116 543454
rect 9352 543218 9436 543454
rect 9672 543218 31258 543454
rect 31494 543218 31578 543454
rect 31814 543218 35617 543454
rect 35853 543218 132653 543454
rect 132889 543218 139589 543454
rect 139825 543218 236625 543454
rect 236861 543218 248858 543454
rect 249094 543218 249178 543454
rect 249414 543218 276058 543454
rect 276294 543218 276378 543454
rect 276614 543218 303258 543454
rect 303494 543218 303578 543454
rect 303814 543218 330458 543454
rect 330694 543218 330778 543454
rect 331014 543218 342545 543454
rect 342781 543218 439581 543454
rect 439817 543218 446517 543454
rect 446753 543218 543553 543454
rect 543789 543218 548058 543454
rect 548294 543218 548378 543454
rect 548614 543218 570292 543454
rect 570528 543218 570612 543454
rect 570848 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 9116 543134
rect 9352 542898 9436 543134
rect 9672 542898 31258 543134
rect 31494 542898 31578 543134
rect 31814 542898 35617 543134
rect 35853 542898 132653 543134
rect 132889 542898 139589 543134
rect 139825 542898 236625 543134
rect 236861 542898 248858 543134
rect 249094 542898 249178 543134
rect 249414 542898 276058 543134
rect 276294 542898 276378 543134
rect 276614 542898 303258 543134
rect 303494 542898 303578 543134
rect 303814 542898 330458 543134
rect 330694 542898 330778 543134
rect 331014 542898 342545 543134
rect 342781 542898 439581 543134
rect 439817 542898 446517 543134
rect 446753 542898 543553 543134
rect 543789 542898 548058 543134
rect 548294 542898 548378 543134
rect 548614 542898 570292 543134
rect 570528 542898 570612 543134
rect 570848 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 7876 525454
rect 8112 525218 8196 525454
rect 8432 525218 17658 525454
rect 17894 525218 17978 525454
rect 18214 525218 44858 525454
rect 45094 525218 45178 525454
rect 45414 525218 72058 525454
rect 72294 525218 72378 525454
rect 72614 525218 99258 525454
rect 99494 525218 99578 525454
rect 99814 525218 126458 525454
rect 126694 525218 126778 525454
rect 127014 525218 153658 525454
rect 153894 525218 153978 525454
rect 154214 525218 180858 525454
rect 181094 525218 181178 525454
rect 181414 525218 208058 525454
rect 208294 525218 208378 525454
rect 208614 525218 235258 525454
rect 235494 525218 235578 525454
rect 235814 525218 262458 525454
rect 262694 525218 262778 525454
rect 263014 525218 289658 525454
rect 289894 525218 289978 525454
rect 290214 525218 316858 525454
rect 317094 525218 317178 525454
rect 317414 525218 344058 525454
rect 344294 525218 344378 525454
rect 344614 525218 371258 525454
rect 371494 525218 371578 525454
rect 371814 525218 398458 525454
rect 398694 525218 398778 525454
rect 399014 525218 425658 525454
rect 425894 525218 425978 525454
rect 426214 525218 452858 525454
rect 453094 525218 453178 525454
rect 453414 525218 480058 525454
rect 480294 525218 480378 525454
rect 480614 525218 507258 525454
rect 507494 525218 507578 525454
rect 507814 525218 534458 525454
rect 534694 525218 534778 525454
rect 535014 525218 561658 525454
rect 561894 525218 561978 525454
rect 562214 525218 571532 525454
rect 571768 525218 571852 525454
rect 572088 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 7876 525134
rect 8112 524898 8196 525134
rect 8432 524898 17658 525134
rect 17894 524898 17978 525134
rect 18214 524898 44858 525134
rect 45094 524898 45178 525134
rect 45414 524898 72058 525134
rect 72294 524898 72378 525134
rect 72614 524898 99258 525134
rect 99494 524898 99578 525134
rect 99814 524898 126458 525134
rect 126694 524898 126778 525134
rect 127014 524898 153658 525134
rect 153894 524898 153978 525134
rect 154214 524898 180858 525134
rect 181094 524898 181178 525134
rect 181414 524898 208058 525134
rect 208294 524898 208378 525134
rect 208614 524898 235258 525134
rect 235494 524898 235578 525134
rect 235814 524898 262458 525134
rect 262694 524898 262778 525134
rect 263014 524898 289658 525134
rect 289894 524898 289978 525134
rect 290214 524898 316858 525134
rect 317094 524898 317178 525134
rect 317414 524898 344058 525134
rect 344294 524898 344378 525134
rect 344614 524898 371258 525134
rect 371494 524898 371578 525134
rect 371814 524898 398458 525134
rect 398694 524898 398778 525134
rect 399014 524898 425658 525134
rect 425894 524898 425978 525134
rect 426214 524898 452858 525134
rect 453094 524898 453178 525134
rect 453414 524898 480058 525134
rect 480294 524898 480378 525134
rect 480614 524898 507258 525134
rect 507494 524898 507578 525134
rect 507814 524898 534458 525134
rect 534694 524898 534778 525134
rect 535014 524898 561658 525134
rect 561894 524898 561978 525134
rect 562214 524898 571532 525134
rect 571768 524898 571852 525134
rect 572088 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 9116 507454
rect 9352 507218 9436 507454
rect 9672 507218 31258 507454
rect 31494 507218 31578 507454
rect 31814 507218 35617 507454
rect 35853 507218 132653 507454
rect 132889 507218 139589 507454
rect 139825 507218 236625 507454
rect 236861 507218 248858 507454
rect 249094 507218 249178 507454
rect 249414 507218 276058 507454
rect 276294 507218 276378 507454
rect 276614 507218 303258 507454
rect 303494 507218 303578 507454
rect 303814 507218 330458 507454
rect 330694 507218 330778 507454
rect 331014 507218 342545 507454
rect 342781 507218 439581 507454
rect 439817 507218 446517 507454
rect 446753 507218 543553 507454
rect 543789 507218 548058 507454
rect 548294 507218 548378 507454
rect 548614 507218 570292 507454
rect 570528 507218 570612 507454
rect 570848 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 9116 507134
rect 9352 506898 9436 507134
rect 9672 506898 31258 507134
rect 31494 506898 31578 507134
rect 31814 506898 35617 507134
rect 35853 506898 132653 507134
rect 132889 506898 139589 507134
rect 139825 506898 236625 507134
rect 236861 506898 248858 507134
rect 249094 506898 249178 507134
rect 249414 506898 276058 507134
rect 276294 506898 276378 507134
rect 276614 506898 303258 507134
rect 303494 506898 303578 507134
rect 303814 506898 330458 507134
rect 330694 506898 330778 507134
rect 331014 506898 342545 507134
rect 342781 506898 439581 507134
rect 439817 506898 446517 507134
rect 446753 506898 543553 507134
rect 543789 506898 548058 507134
rect 548294 506898 548378 507134
rect 548614 506898 570292 507134
rect 570528 506898 570612 507134
rect 570848 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 7876 489454
rect 8112 489218 8196 489454
rect 8432 489218 17658 489454
rect 17894 489218 17978 489454
rect 18214 489218 34897 489454
rect 35133 489218 133373 489454
rect 133609 489218 138869 489454
rect 139105 489218 237345 489454
rect 237581 489218 262458 489454
rect 262694 489218 262778 489454
rect 263014 489218 289658 489454
rect 289894 489218 289978 489454
rect 290214 489218 316858 489454
rect 317094 489218 317178 489454
rect 317414 489218 341825 489454
rect 342061 489218 440301 489454
rect 440537 489218 445797 489454
rect 446033 489218 544273 489454
rect 544509 489218 561658 489454
rect 561894 489218 561978 489454
rect 562214 489218 571532 489454
rect 571768 489218 571852 489454
rect 572088 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 7876 489134
rect 8112 488898 8196 489134
rect 8432 488898 17658 489134
rect 17894 488898 17978 489134
rect 18214 488898 34897 489134
rect 35133 488898 133373 489134
rect 133609 488898 138869 489134
rect 139105 488898 237345 489134
rect 237581 488898 262458 489134
rect 262694 488898 262778 489134
rect 263014 488898 289658 489134
rect 289894 488898 289978 489134
rect 290214 488898 316858 489134
rect 317094 488898 317178 489134
rect 317414 488898 341825 489134
rect 342061 488898 440301 489134
rect 440537 488898 445797 489134
rect 446033 488898 544273 489134
rect 544509 488898 561658 489134
rect 561894 488898 561978 489134
rect 562214 488898 571532 489134
rect 571768 488898 571852 489134
rect 572088 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 9116 471454
rect 9352 471218 9436 471454
rect 9672 471218 31258 471454
rect 31494 471218 31578 471454
rect 31814 471218 35617 471454
rect 35853 471218 132653 471454
rect 132889 471218 139589 471454
rect 139825 471218 236625 471454
rect 236861 471218 248858 471454
rect 249094 471218 249178 471454
rect 249414 471218 276058 471454
rect 276294 471218 276378 471454
rect 276614 471218 303258 471454
rect 303494 471218 303578 471454
rect 303814 471218 330458 471454
rect 330694 471218 330778 471454
rect 331014 471218 342545 471454
rect 342781 471218 439581 471454
rect 439817 471218 446517 471454
rect 446753 471218 543553 471454
rect 543789 471218 548058 471454
rect 548294 471218 548378 471454
rect 548614 471218 570292 471454
rect 570528 471218 570612 471454
rect 570848 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 9116 471134
rect 9352 470898 9436 471134
rect 9672 470898 31258 471134
rect 31494 470898 31578 471134
rect 31814 470898 35617 471134
rect 35853 470898 132653 471134
rect 132889 470898 139589 471134
rect 139825 470898 236625 471134
rect 236861 470898 248858 471134
rect 249094 470898 249178 471134
rect 249414 470898 276058 471134
rect 276294 470898 276378 471134
rect 276614 470898 303258 471134
rect 303494 470898 303578 471134
rect 303814 470898 330458 471134
rect 330694 470898 330778 471134
rect 331014 470898 342545 471134
rect 342781 470898 439581 471134
rect 439817 470898 446517 471134
rect 446753 470898 543553 471134
rect 543789 470898 548058 471134
rect 548294 470898 548378 471134
rect 548614 470898 570292 471134
rect 570528 470898 570612 471134
rect 570848 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 7876 453454
rect 8112 453218 8196 453454
rect 8432 453218 17658 453454
rect 17894 453218 17978 453454
rect 18214 453218 34897 453454
rect 35133 453218 133373 453454
rect 133609 453218 138869 453454
rect 139105 453218 237345 453454
rect 237581 453218 262458 453454
rect 262694 453218 262778 453454
rect 263014 453218 289658 453454
rect 289894 453218 289978 453454
rect 290214 453218 316858 453454
rect 317094 453218 317178 453454
rect 317414 453218 341825 453454
rect 342061 453218 440301 453454
rect 440537 453218 445797 453454
rect 446033 453218 544273 453454
rect 544509 453218 561658 453454
rect 561894 453218 561978 453454
rect 562214 453218 571532 453454
rect 571768 453218 571852 453454
rect 572088 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 7876 453134
rect 8112 452898 8196 453134
rect 8432 452898 17658 453134
rect 17894 452898 17978 453134
rect 18214 452898 34897 453134
rect 35133 452898 133373 453134
rect 133609 452898 138869 453134
rect 139105 452898 237345 453134
rect 237581 452898 262458 453134
rect 262694 452898 262778 453134
rect 263014 452898 289658 453134
rect 289894 452898 289978 453134
rect 290214 452898 316858 453134
rect 317094 452898 317178 453134
rect 317414 452898 341825 453134
rect 342061 452898 440301 453134
rect 440537 452898 445797 453134
rect 446033 452898 544273 453134
rect 544509 452898 561658 453134
rect 561894 452898 561978 453134
rect 562214 452898 571532 453134
rect 571768 452898 571852 453134
rect 572088 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 9116 435454
rect 9352 435218 9436 435454
rect 9672 435218 31258 435454
rect 31494 435218 31578 435454
rect 31814 435218 58458 435454
rect 58694 435218 58778 435454
rect 59014 435218 85658 435454
rect 85894 435218 85978 435454
rect 86214 435218 112858 435454
rect 113094 435218 113178 435454
rect 113414 435218 140058 435454
rect 140294 435218 140378 435454
rect 140614 435218 167258 435454
rect 167494 435218 167578 435454
rect 167814 435218 194458 435454
rect 194694 435218 194778 435454
rect 195014 435218 221658 435454
rect 221894 435218 221978 435454
rect 222214 435218 248858 435454
rect 249094 435218 249178 435454
rect 249414 435218 276058 435454
rect 276294 435218 276378 435454
rect 276614 435218 303258 435454
rect 303494 435218 303578 435454
rect 303814 435218 330458 435454
rect 330694 435218 330778 435454
rect 331014 435218 357658 435454
rect 357894 435218 357978 435454
rect 358214 435218 384858 435454
rect 385094 435218 385178 435454
rect 385414 435218 412058 435454
rect 412294 435218 412378 435454
rect 412614 435218 439258 435454
rect 439494 435218 439578 435454
rect 439814 435218 466458 435454
rect 466694 435218 466778 435454
rect 467014 435218 493658 435454
rect 493894 435218 493978 435454
rect 494214 435218 520858 435454
rect 521094 435218 521178 435454
rect 521414 435218 548058 435454
rect 548294 435218 548378 435454
rect 548614 435218 570292 435454
rect 570528 435218 570612 435454
rect 570848 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 9116 435134
rect 9352 434898 9436 435134
rect 9672 434898 31258 435134
rect 31494 434898 31578 435134
rect 31814 434898 58458 435134
rect 58694 434898 58778 435134
rect 59014 434898 85658 435134
rect 85894 434898 85978 435134
rect 86214 434898 112858 435134
rect 113094 434898 113178 435134
rect 113414 434898 140058 435134
rect 140294 434898 140378 435134
rect 140614 434898 167258 435134
rect 167494 434898 167578 435134
rect 167814 434898 194458 435134
rect 194694 434898 194778 435134
rect 195014 434898 221658 435134
rect 221894 434898 221978 435134
rect 222214 434898 248858 435134
rect 249094 434898 249178 435134
rect 249414 434898 276058 435134
rect 276294 434898 276378 435134
rect 276614 434898 303258 435134
rect 303494 434898 303578 435134
rect 303814 434898 330458 435134
rect 330694 434898 330778 435134
rect 331014 434898 357658 435134
rect 357894 434898 357978 435134
rect 358214 434898 384858 435134
rect 385094 434898 385178 435134
rect 385414 434898 412058 435134
rect 412294 434898 412378 435134
rect 412614 434898 439258 435134
rect 439494 434898 439578 435134
rect 439814 434898 466458 435134
rect 466694 434898 466778 435134
rect 467014 434898 493658 435134
rect 493894 434898 493978 435134
rect 494214 434898 520858 435134
rect 521094 434898 521178 435134
rect 521414 434898 548058 435134
rect 548294 434898 548378 435134
rect 548614 434898 570292 435134
rect 570528 434898 570612 435134
rect 570848 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 7876 417454
rect 8112 417218 8196 417454
rect 8432 417218 17658 417454
rect 17894 417218 17978 417454
rect 18214 417218 44858 417454
rect 45094 417218 45178 417454
rect 45414 417218 72058 417454
rect 72294 417218 72378 417454
rect 72614 417218 99258 417454
rect 99494 417218 99578 417454
rect 99814 417218 126458 417454
rect 126694 417218 126778 417454
rect 127014 417218 153658 417454
rect 153894 417218 153978 417454
rect 154214 417218 180858 417454
rect 181094 417218 181178 417454
rect 181414 417218 208058 417454
rect 208294 417218 208378 417454
rect 208614 417218 235258 417454
rect 235494 417218 235578 417454
rect 235814 417218 262458 417454
rect 262694 417218 262778 417454
rect 263014 417218 289658 417454
rect 289894 417218 289978 417454
rect 290214 417218 316858 417454
rect 317094 417218 317178 417454
rect 317414 417218 341825 417454
rect 342061 417218 440301 417454
rect 440537 417218 445797 417454
rect 446033 417218 544273 417454
rect 544509 417218 561658 417454
rect 561894 417218 561978 417454
rect 562214 417218 571532 417454
rect 571768 417218 571852 417454
rect 572088 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 7876 417134
rect 8112 416898 8196 417134
rect 8432 416898 17658 417134
rect 17894 416898 17978 417134
rect 18214 416898 44858 417134
rect 45094 416898 45178 417134
rect 45414 416898 72058 417134
rect 72294 416898 72378 417134
rect 72614 416898 99258 417134
rect 99494 416898 99578 417134
rect 99814 416898 126458 417134
rect 126694 416898 126778 417134
rect 127014 416898 153658 417134
rect 153894 416898 153978 417134
rect 154214 416898 180858 417134
rect 181094 416898 181178 417134
rect 181414 416898 208058 417134
rect 208294 416898 208378 417134
rect 208614 416898 235258 417134
rect 235494 416898 235578 417134
rect 235814 416898 262458 417134
rect 262694 416898 262778 417134
rect 263014 416898 289658 417134
rect 289894 416898 289978 417134
rect 290214 416898 316858 417134
rect 317094 416898 317178 417134
rect 317414 416898 341825 417134
rect 342061 416898 440301 417134
rect 440537 416898 445797 417134
rect 446033 416898 544273 417134
rect 544509 416898 561658 417134
rect 561894 416898 561978 417134
rect 562214 416898 571532 417134
rect 571768 416898 571852 417134
rect 572088 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 9116 399454
rect 9352 399218 9436 399454
rect 9672 399218 31258 399454
rect 31494 399218 31578 399454
rect 31814 399218 58458 399454
rect 58694 399218 58778 399454
rect 59014 399218 85658 399454
rect 85894 399218 85978 399454
rect 86214 399218 112858 399454
rect 113094 399218 113178 399454
rect 113414 399218 140058 399454
rect 140294 399218 140378 399454
rect 140614 399218 167258 399454
rect 167494 399218 167578 399454
rect 167814 399218 194458 399454
rect 194694 399218 194778 399454
rect 195014 399218 221658 399454
rect 221894 399218 221978 399454
rect 222214 399218 248858 399454
rect 249094 399218 249178 399454
rect 249414 399218 276058 399454
rect 276294 399218 276378 399454
rect 276614 399218 303258 399454
rect 303494 399218 303578 399454
rect 303814 399218 330458 399454
rect 330694 399218 330778 399454
rect 331014 399218 342545 399454
rect 342781 399218 439581 399454
rect 439817 399218 446517 399454
rect 446753 399218 543553 399454
rect 543789 399218 548058 399454
rect 548294 399218 548378 399454
rect 548614 399218 570292 399454
rect 570528 399218 570612 399454
rect 570848 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 9116 399134
rect 9352 398898 9436 399134
rect 9672 398898 31258 399134
rect 31494 398898 31578 399134
rect 31814 398898 58458 399134
rect 58694 398898 58778 399134
rect 59014 398898 85658 399134
rect 85894 398898 85978 399134
rect 86214 398898 112858 399134
rect 113094 398898 113178 399134
rect 113414 398898 140058 399134
rect 140294 398898 140378 399134
rect 140614 398898 167258 399134
rect 167494 398898 167578 399134
rect 167814 398898 194458 399134
rect 194694 398898 194778 399134
rect 195014 398898 221658 399134
rect 221894 398898 221978 399134
rect 222214 398898 248858 399134
rect 249094 398898 249178 399134
rect 249414 398898 276058 399134
rect 276294 398898 276378 399134
rect 276614 398898 303258 399134
rect 303494 398898 303578 399134
rect 303814 398898 330458 399134
rect 330694 398898 330778 399134
rect 331014 398898 342545 399134
rect 342781 398898 439581 399134
rect 439817 398898 446517 399134
rect 446753 398898 543553 399134
rect 543789 398898 548058 399134
rect 548294 398898 548378 399134
rect 548614 398898 570292 399134
rect 570528 398898 570612 399134
rect 570848 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 7876 381454
rect 8112 381218 8196 381454
rect 8432 381218 17658 381454
rect 17894 381218 17978 381454
rect 18214 381218 44858 381454
rect 45094 381218 45178 381454
rect 45414 381218 72058 381454
rect 72294 381218 72378 381454
rect 72614 381218 99258 381454
rect 99494 381218 99578 381454
rect 99814 381218 126458 381454
rect 126694 381218 126778 381454
rect 127014 381218 153658 381454
rect 153894 381218 153978 381454
rect 154214 381218 180858 381454
rect 181094 381218 181178 381454
rect 181414 381218 208058 381454
rect 208294 381218 208378 381454
rect 208614 381218 235258 381454
rect 235494 381218 235578 381454
rect 235814 381218 262458 381454
rect 262694 381218 262778 381454
rect 263014 381218 289658 381454
rect 289894 381218 289978 381454
rect 290214 381218 316858 381454
rect 317094 381218 317178 381454
rect 317414 381218 341825 381454
rect 342061 381218 440301 381454
rect 440537 381218 445797 381454
rect 446033 381218 544273 381454
rect 544509 381218 561658 381454
rect 561894 381218 561978 381454
rect 562214 381218 571532 381454
rect 571768 381218 571852 381454
rect 572088 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 7876 381134
rect 8112 380898 8196 381134
rect 8432 380898 17658 381134
rect 17894 380898 17978 381134
rect 18214 380898 44858 381134
rect 45094 380898 45178 381134
rect 45414 380898 72058 381134
rect 72294 380898 72378 381134
rect 72614 380898 99258 381134
rect 99494 380898 99578 381134
rect 99814 380898 126458 381134
rect 126694 380898 126778 381134
rect 127014 380898 153658 381134
rect 153894 380898 153978 381134
rect 154214 380898 180858 381134
rect 181094 380898 181178 381134
rect 181414 380898 208058 381134
rect 208294 380898 208378 381134
rect 208614 380898 235258 381134
rect 235494 380898 235578 381134
rect 235814 380898 262458 381134
rect 262694 380898 262778 381134
rect 263014 380898 289658 381134
rect 289894 380898 289978 381134
rect 290214 380898 316858 381134
rect 317094 380898 317178 381134
rect 317414 380898 341825 381134
rect 342061 380898 440301 381134
rect 440537 380898 445797 381134
rect 446033 380898 544273 381134
rect 544509 380898 561658 381134
rect 561894 380898 561978 381134
rect 562214 380898 571532 381134
rect 571768 380898 571852 381134
rect 572088 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 9116 363454
rect 9352 363218 9436 363454
rect 9672 363218 31258 363454
rect 31494 363218 31578 363454
rect 31814 363218 35617 363454
rect 35853 363218 132653 363454
rect 132889 363218 139589 363454
rect 139825 363218 236625 363454
rect 236861 363218 248858 363454
rect 249094 363218 249178 363454
rect 249414 363218 276058 363454
rect 276294 363218 276378 363454
rect 276614 363218 303258 363454
rect 303494 363218 303578 363454
rect 303814 363218 330458 363454
rect 330694 363218 330778 363454
rect 331014 363218 342545 363454
rect 342781 363218 439581 363454
rect 439817 363218 446517 363454
rect 446753 363218 543553 363454
rect 543789 363218 548058 363454
rect 548294 363218 548378 363454
rect 548614 363218 570292 363454
rect 570528 363218 570612 363454
rect 570848 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 9116 363134
rect 9352 362898 9436 363134
rect 9672 362898 31258 363134
rect 31494 362898 31578 363134
rect 31814 362898 35617 363134
rect 35853 362898 132653 363134
rect 132889 362898 139589 363134
rect 139825 362898 236625 363134
rect 236861 362898 248858 363134
rect 249094 362898 249178 363134
rect 249414 362898 276058 363134
rect 276294 362898 276378 363134
rect 276614 362898 303258 363134
rect 303494 362898 303578 363134
rect 303814 362898 330458 363134
rect 330694 362898 330778 363134
rect 331014 362898 342545 363134
rect 342781 362898 439581 363134
rect 439817 362898 446517 363134
rect 446753 362898 543553 363134
rect 543789 362898 548058 363134
rect 548294 362898 548378 363134
rect 548614 362898 570292 363134
rect 570528 362898 570612 363134
rect 570848 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 7876 345454
rect 8112 345218 8196 345454
rect 8432 345218 17658 345454
rect 17894 345218 17978 345454
rect 18214 345218 34897 345454
rect 35133 345218 133373 345454
rect 133609 345218 138869 345454
rect 139105 345218 237345 345454
rect 237581 345218 262458 345454
rect 262694 345218 262778 345454
rect 263014 345218 289658 345454
rect 289894 345218 289978 345454
rect 290214 345218 316858 345454
rect 317094 345218 317178 345454
rect 317414 345218 341825 345454
rect 342061 345218 440301 345454
rect 440537 345218 445797 345454
rect 446033 345218 544273 345454
rect 544509 345218 561658 345454
rect 561894 345218 561978 345454
rect 562214 345218 571532 345454
rect 571768 345218 571852 345454
rect 572088 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 7876 345134
rect 8112 344898 8196 345134
rect 8432 344898 17658 345134
rect 17894 344898 17978 345134
rect 18214 344898 34897 345134
rect 35133 344898 133373 345134
rect 133609 344898 138869 345134
rect 139105 344898 237345 345134
rect 237581 344898 262458 345134
rect 262694 344898 262778 345134
rect 263014 344898 289658 345134
rect 289894 344898 289978 345134
rect 290214 344898 316858 345134
rect 317094 344898 317178 345134
rect 317414 344898 341825 345134
rect 342061 344898 440301 345134
rect 440537 344898 445797 345134
rect 446033 344898 544273 345134
rect 544509 344898 561658 345134
rect 561894 344898 561978 345134
rect 562214 344898 571532 345134
rect 571768 344898 571852 345134
rect 572088 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 9116 327454
rect 9352 327218 9436 327454
rect 9672 327218 31258 327454
rect 31494 327218 31578 327454
rect 31814 327218 35617 327454
rect 35853 327218 132653 327454
rect 132889 327218 139589 327454
rect 139825 327218 236625 327454
rect 236861 327218 248858 327454
rect 249094 327218 249178 327454
rect 249414 327218 276058 327454
rect 276294 327218 276378 327454
rect 276614 327218 303258 327454
rect 303494 327218 303578 327454
rect 303814 327218 330458 327454
rect 330694 327218 330778 327454
rect 331014 327218 342545 327454
rect 342781 327218 446517 327454
rect 446753 327218 543553 327454
rect 543789 327218 548058 327454
rect 548294 327218 548378 327454
rect 548614 327218 570292 327454
rect 570528 327218 570612 327454
rect 570848 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 9116 327134
rect 9352 326898 9436 327134
rect 9672 326898 31258 327134
rect 31494 326898 31578 327134
rect 31814 326898 35617 327134
rect 35853 326898 132653 327134
rect 132889 326898 139589 327134
rect 139825 326898 236625 327134
rect 236861 326898 248858 327134
rect 249094 326898 249178 327134
rect 249414 326898 276058 327134
rect 276294 326898 276378 327134
rect 276614 326898 303258 327134
rect 303494 326898 303578 327134
rect 303814 326898 330458 327134
rect 330694 326898 330778 327134
rect 331014 326898 342545 327134
rect 342781 326898 446517 327134
rect 446753 326898 543553 327134
rect 543789 326898 548058 327134
rect 548294 326898 548378 327134
rect 548614 326898 570292 327134
rect 570528 326898 570612 327134
rect 570848 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 7876 309454
rect 8112 309218 8196 309454
rect 8432 309218 17658 309454
rect 17894 309218 17978 309454
rect 18214 309218 34897 309454
rect 35133 309218 133373 309454
rect 133609 309218 138869 309454
rect 139105 309218 237345 309454
rect 237581 309218 262458 309454
rect 262694 309218 262778 309454
rect 263014 309218 289658 309454
rect 289894 309218 289978 309454
rect 290214 309218 316858 309454
rect 317094 309218 317178 309454
rect 317414 309218 341825 309454
rect 342061 309218 440301 309454
rect 440537 309218 445797 309454
rect 446033 309218 544273 309454
rect 544509 309218 561658 309454
rect 561894 309218 561978 309454
rect 562214 309218 571532 309454
rect 571768 309218 571852 309454
rect 572088 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 7876 309134
rect 8112 308898 8196 309134
rect 8432 308898 17658 309134
rect 17894 308898 17978 309134
rect 18214 308898 34897 309134
rect 35133 308898 133373 309134
rect 133609 308898 138869 309134
rect 139105 308898 237345 309134
rect 237581 308898 262458 309134
rect 262694 308898 262778 309134
rect 263014 308898 289658 309134
rect 289894 308898 289978 309134
rect 290214 308898 316858 309134
rect 317094 308898 317178 309134
rect 317414 308898 341825 309134
rect 342061 308898 440301 309134
rect 440537 308898 445797 309134
rect 446033 308898 544273 309134
rect 544509 308898 561658 309134
rect 561894 308898 561978 309134
rect 562214 308898 571532 309134
rect 571768 308898 571852 309134
rect 572088 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 9116 291454
rect 9352 291218 9436 291454
rect 9672 291218 31258 291454
rect 31494 291218 31578 291454
rect 31814 291218 35617 291454
rect 35853 291218 132653 291454
rect 132889 291218 139589 291454
rect 139825 291218 236625 291454
rect 236861 291218 248858 291454
rect 249094 291218 249178 291454
rect 249414 291218 276058 291454
rect 276294 291218 276378 291454
rect 276614 291218 303258 291454
rect 303494 291218 303578 291454
rect 303814 291218 330458 291454
rect 330694 291218 330778 291454
rect 331014 291218 342545 291454
rect 342781 291218 439581 291454
rect 439817 291218 446517 291454
rect 446753 291218 543553 291454
rect 543789 291218 548058 291454
rect 548294 291218 548378 291454
rect 548614 291218 570292 291454
rect 570528 291218 570612 291454
rect 570848 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 9116 291134
rect 9352 290898 9436 291134
rect 9672 290898 31258 291134
rect 31494 290898 31578 291134
rect 31814 290898 35617 291134
rect 35853 290898 132653 291134
rect 132889 290898 139589 291134
rect 139825 290898 236625 291134
rect 236861 290898 248858 291134
rect 249094 290898 249178 291134
rect 249414 290898 276058 291134
rect 276294 290898 276378 291134
rect 276614 290898 303258 291134
rect 303494 290898 303578 291134
rect 303814 290898 330458 291134
rect 330694 290898 330778 291134
rect 331014 290898 342545 291134
rect 342781 290898 439581 291134
rect 439817 290898 446517 291134
rect 446753 290898 543553 291134
rect 543789 290898 548058 291134
rect 548294 290898 548378 291134
rect 548614 290898 570292 291134
rect 570528 290898 570612 291134
rect 570848 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 7876 273454
rect 8112 273218 8196 273454
rect 8432 273218 17658 273454
rect 17894 273218 17978 273454
rect 18214 273218 44858 273454
rect 45094 273218 45178 273454
rect 45414 273218 72058 273454
rect 72294 273218 72378 273454
rect 72614 273218 99258 273454
rect 99494 273218 99578 273454
rect 99814 273218 126458 273454
rect 126694 273218 126778 273454
rect 127014 273218 153658 273454
rect 153894 273218 153978 273454
rect 154214 273218 180858 273454
rect 181094 273218 181178 273454
rect 181414 273218 208058 273454
rect 208294 273218 208378 273454
rect 208614 273218 235258 273454
rect 235494 273218 235578 273454
rect 235814 273218 262458 273454
rect 262694 273218 262778 273454
rect 263014 273218 289658 273454
rect 289894 273218 289978 273454
rect 290214 273218 316858 273454
rect 317094 273218 317178 273454
rect 317414 273218 341825 273454
rect 342061 273218 440301 273454
rect 440537 273218 445797 273454
rect 446033 273218 544273 273454
rect 544509 273218 561658 273454
rect 561894 273218 561978 273454
rect 562214 273218 571532 273454
rect 571768 273218 571852 273454
rect 572088 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 7876 273134
rect 8112 272898 8196 273134
rect 8432 272898 17658 273134
rect 17894 272898 17978 273134
rect 18214 272898 44858 273134
rect 45094 272898 45178 273134
rect 45414 272898 72058 273134
rect 72294 272898 72378 273134
rect 72614 272898 99258 273134
rect 99494 272898 99578 273134
rect 99814 272898 126458 273134
rect 126694 272898 126778 273134
rect 127014 272898 153658 273134
rect 153894 272898 153978 273134
rect 154214 272898 180858 273134
rect 181094 272898 181178 273134
rect 181414 272898 208058 273134
rect 208294 272898 208378 273134
rect 208614 272898 235258 273134
rect 235494 272898 235578 273134
rect 235814 272898 262458 273134
rect 262694 272898 262778 273134
rect 263014 272898 289658 273134
rect 289894 272898 289978 273134
rect 290214 272898 316858 273134
rect 317094 272898 317178 273134
rect 317414 272898 341825 273134
rect 342061 272898 440301 273134
rect 440537 272898 445797 273134
rect 446033 272898 544273 273134
rect 544509 272898 561658 273134
rect 561894 272898 561978 273134
rect 562214 272898 571532 273134
rect 571768 272898 571852 273134
rect 572088 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 9116 255454
rect 9352 255218 9436 255454
rect 9672 255218 31258 255454
rect 31494 255218 31578 255454
rect 31814 255218 58458 255454
rect 58694 255218 58778 255454
rect 59014 255218 85658 255454
rect 85894 255218 85978 255454
rect 86214 255218 112858 255454
rect 113094 255218 113178 255454
rect 113414 255218 140058 255454
rect 140294 255218 140378 255454
rect 140614 255218 167258 255454
rect 167494 255218 167578 255454
rect 167814 255218 194458 255454
rect 194694 255218 194778 255454
rect 195014 255218 221658 255454
rect 221894 255218 221978 255454
rect 222214 255218 248858 255454
rect 249094 255218 249178 255454
rect 249414 255218 276058 255454
rect 276294 255218 276378 255454
rect 276614 255218 303258 255454
rect 303494 255218 303578 255454
rect 303814 255218 330458 255454
rect 330694 255218 330778 255454
rect 331014 255218 342545 255454
rect 342781 255218 439581 255454
rect 439817 255218 446517 255454
rect 446753 255218 543553 255454
rect 543789 255218 548058 255454
rect 548294 255218 548378 255454
rect 548614 255218 570292 255454
rect 570528 255218 570612 255454
rect 570848 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 9116 255134
rect 9352 254898 9436 255134
rect 9672 254898 31258 255134
rect 31494 254898 31578 255134
rect 31814 254898 58458 255134
rect 58694 254898 58778 255134
rect 59014 254898 85658 255134
rect 85894 254898 85978 255134
rect 86214 254898 112858 255134
rect 113094 254898 113178 255134
rect 113414 254898 140058 255134
rect 140294 254898 140378 255134
rect 140614 254898 167258 255134
rect 167494 254898 167578 255134
rect 167814 254898 194458 255134
rect 194694 254898 194778 255134
rect 195014 254898 221658 255134
rect 221894 254898 221978 255134
rect 222214 254898 248858 255134
rect 249094 254898 249178 255134
rect 249414 254898 276058 255134
rect 276294 254898 276378 255134
rect 276614 254898 303258 255134
rect 303494 254898 303578 255134
rect 303814 254898 330458 255134
rect 330694 254898 330778 255134
rect 331014 254898 342545 255134
rect 342781 254898 439581 255134
rect 439817 254898 446517 255134
rect 446753 254898 543553 255134
rect 543789 254898 548058 255134
rect 548294 254898 548378 255134
rect 548614 254898 570292 255134
rect 570528 254898 570612 255134
rect 570848 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 7876 237454
rect 8112 237218 8196 237454
rect 8432 237218 17658 237454
rect 17894 237218 17978 237454
rect 18214 237218 44858 237454
rect 45094 237218 45178 237454
rect 45414 237218 72058 237454
rect 72294 237218 72378 237454
rect 72614 237218 99258 237454
rect 99494 237218 99578 237454
rect 99814 237218 126458 237454
rect 126694 237218 126778 237454
rect 127014 237218 153658 237454
rect 153894 237218 153978 237454
rect 154214 237218 180858 237454
rect 181094 237218 181178 237454
rect 181414 237218 208058 237454
rect 208294 237218 208378 237454
rect 208614 237218 235258 237454
rect 235494 237218 235578 237454
rect 235814 237218 262458 237454
rect 262694 237218 262778 237454
rect 263014 237218 289658 237454
rect 289894 237218 289978 237454
rect 290214 237218 316858 237454
rect 317094 237218 317178 237454
rect 317414 237218 344058 237454
rect 344294 237218 344378 237454
rect 344614 237218 371258 237454
rect 371494 237218 371578 237454
rect 371814 237218 398458 237454
rect 398694 237218 398778 237454
rect 399014 237218 425658 237454
rect 425894 237218 425978 237454
rect 426214 237218 452858 237454
rect 453094 237218 453178 237454
rect 453414 237218 480058 237454
rect 480294 237218 480378 237454
rect 480614 237218 507258 237454
rect 507494 237218 507578 237454
rect 507814 237218 534458 237454
rect 534694 237218 534778 237454
rect 535014 237218 561658 237454
rect 561894 237218 561978 237454
rect 562214 237218 571532 237454
rect 571768 237218 571852 237454
rect 572088 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 7876 237134
rect 8112 236898 8196 237134
rect 8432 236898 17658 237134
rect 17894 236898 17978 237134
rect 18214 236898 44858 237134
rect 45094 236898 45178 237134
rect 45414 236898 72058 237134
rect 72294 236898 72378 237134
rect 72614 236898 99258 237134
rect 99494 236898 99578 237134
rect 99814 236898 126458 237134
rect 126694 236898 126778 237134
rect 127014 236898 153658 237134
rect 153894 236898 153978 237134
rect 154214 236898 180858 237134
rect 181094 236898 181178 237134
rect 181414 236898 208058 237134
rect 208294 236898 208378 237134
rect 208614 236898 235258 237134
rect 235494 236898 235578 237134
rect 235814 236898 262458 237134
rect 262694 236898 262778 237134
rect 263014 236898 289658 237134
rect 289894 236898 289978 237134
rect 290214 236898 316858 237134
rect 317094 236898 317178 237134
rect 317414 236898 344058 237134
rect 344294 236898 344378 237134
rect 344614 236898 371258 237134
rect 371494 236898 371578 237134
rect 371814 236898 398458 237134
rect 398694 236898 398778 237134
rect 399014 236898 425658 237134
rect 425894 236898 425978 237134
rect 426214 236898 452858 237134
rect 453094 236898 453178 237134
rect 453414 236898 480058 237134
rect 480294 236898 480378 237134
rect 480614 236898 507258 237134
rect 507494 236898 507578 237134
rect 507814 236898 534458 237134
rect 534694 236898 534778 237134
rect 535014 236898 561658 237134
rect 561894 236898 561978 237134
rect 562214 236898 571532 237134
rect 571768 236898 571852 237134
rect 572088 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 9116 219454
rect 9352 219218 9436 219454
rect 9672 219218 31258 219454
rect 31494 219218 31578 219454
rect 31814 219218 35617 219454
rect 35853 219218 132653 219454
rect 132889 219218 139589 219454
rect 139825 219218 236625 219454
rect 236861 219218 248858 219454
rect 249094 219218 249178 219454
rect 249414 219218 276058 219454
rect 276294 219218 276378 219454
rect 276614 219218 303258 219454
rect 303494 219218 303578 219454
rect 303814 219218 330458 219454
rect 330694 219218 330778 219454
rect 331014 219218 342545 219454
rect 342781 219218 439581 219454
rect 439817 219218 446517 219454
rect 446753 219218 543553 219454
rect 543789 219218 548058 219454
rect 548294 219218 548378 219454
rect 548614 219218 570292 219454
rect 570528 219218 570612 219454
rect 570848 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 9116 219134
rect 9352 218898 9436 219134
rect 9672 218898 31258 219134
rect 31494 218898 31578 219134
rect 31814 218898 35617 219134
rect 35853 218898 132653 219134
rect 132889 218898 139589 219134
rect 139825 218898 236625 219134
rect 236861 218898 248858 219134
rect 249094 218898 249178 219134
rect 249414 218898 276058 219134
rect 276294 218898 276378 219134
rect 276614 218898 303258 219134
rect 303494 218898 303578 219134
rect 303814 218898 330458 219134
rect 330694 218898 330778 219134
rect 331014 218898 342545 219134
rect 342781 218898 439581 219134
rect 439817 218898 446517 219134
rect 446753 218898 543553 219134
rect 543789 218898 548058 219134
rect 548294 218898 548378 219134
rect 548614 218898 570292 219134
rect 570528 218898 570612 219134
rect 570848 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 7876 201454
rect 8112 201218 8196 201454
rect 8432 201218 17658 201454
rect 17894 201218 17978 201454
rect 18214 201218 34897 201454
rect 35133 201218 133373 201454
rect 133609 201218 138869 201454
rect 139105 201218 237345 201454
rect 237581 201218 262458 201454
rect 262694 201218 262778 201454
rect 263014 201218 289658 201454
rect 289894 201218 289978 201454
rect 290214 201218 316858 201454
rect 317094 201218 317178 201454
rect 317414 201218 341825 201454
rect 342061 201218 440301 201454
rect 440537 201218 445797 201454
rect 446033 201218 544273 201454
rect 544509 201218 561658 201454
rect 561894 201218 561978 201454
rect 562214 201218 571532 201454
rect 571768 201218 571852 201454
rect 572088 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 7876 201134
rect 8112 200898 8196 201134
rect 8432 200898 17658 201134
rect 17894 200898 17978 201134
rect 18214 200898 34897 201134
rect 35133 200898 133373 201134
rect 133609 200898 138869 201134
rect 139105 200898 237345 201134
rect 237581 200898 262458 201134
rect 262694 200898 262778 201134
rect 263014 200898 289658 201134
rect 289894 200898 289978 201134
rect 290214 200898 316858 201134
rect 317094 200898 317178 201134
rect 317414 200898 341825 201134
rect 342061 200898 440301 201134
rect 440537 200898 445797 201134
rect 446033 200898 544273 201134
rect 544509 200898 561658 201134
rect 561894 200898 561978 201134
rect 562214 200898 571532 201134
rect 571768 200898 571852 201134
rect 572088 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 9116 183454
rect 9352 183218 9436 183454
rect 9672 183218 31258 183454
rect 31494 183218 31578 183454
rect 31814 183218 35617 183454
rect 35853 183218 132653 183454
rect 132889 183218 139589 183454
rect 139825 183218 236625 183454
rect 236861 183218 248858 183454
rect 249094 183218 249178 183454
rect 249414 183218 276058 183454
rect 276294 183218 276378 183454
rect 276614 183218 303258 183454
rect 303494 183218 303578 183454
rect 303814 183218 330458 183454
rect 330694 183218 330778 183454
rect 331014 183218 342545 183454
rect 342781 183218 439581 183454
rect 439817 183218 446517 183454
rect 446753 183218 543553 183454
rect 543789 183218 548058 183454
rect 548294 183218 548378 183454
rect 548614 183218 570292 183454
rect 570528 183218 570612 183454
rect 570848 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 9116 183134
rect 9352 182898 9436 183134
rect 9672 182898 31258 183134
rect 31494 182898 31578 183134
rect 31814 182898 35617 183134
rect 35853 182898 132653 183134
rect 132889 182898 139589 183134
rect 139825 182898 236625 183134
rect 236861 182898 248858 183134
rect 249094 182898 249178 183134
rect 249414 182898 276058 183134
rect 276294 182898 276378 183134
rect 276614 182898 303258 183134
rect 303494 182898 303578 183134
rect 303814 182898 330458 183134
rect 330694 182898 330778 183134
rect 331014 182898 342545 183134
rect 342781 182898 439581 183134
rect 439817 182898 446517 183134
rect 446753 182898 543553 183134
rect 543789 182898 548058 183134
rect 548294 182898 548378 183134
rect 548614 182898 570292 183134
rect 570528 182898 570612 183134
rect 570848 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 7876 165454
rect 8112 165218 8196 165454
rect 8432 165218 17658 165454
rect 17894 165218 17978 165454
rect 18214 165218 34897 165454
rect 35133 165218 133373 165454
rect 133609 165218 138869 165454
rect 139105 165218 237345 165454
rect 237581 165218 262458 165454
rect 262694 165218 262778 165454
rect 263014 165218 289658 165454
rect 289894 165218 289978 165454
rect 290214 165218 316858 165454
rect 317094 165218 317178 165454
rect 317414 165218 341825 165454
rect 342061 165218 440301 165454
rect 440537 165218 445797 165454
rect 446033 165218 544273 165454
rect 544509 165218 561658 165454
rect 561894 165218 561978 165454
rect 562214 165218 571532 165454
rect 571768 165218 571852 165454
rect 572088 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 7876 165134
rect 8112 164898 8196 165134
rect 8432 164898 17658 165134
rect 17894 164898 17978 165134
rect 18214 164898 34897 165134
rect 35133 164898 133373 165134
rect 133609 164898 138869 165134
rect 139105 164898 237345 165134
rect 237581 164898 262458 165134
rect 262694 164898 262778 165134
rect 263014 164898 289658 165134
rect 289894 164898 289978 165134
rect 290214 164898 316858 165134
rect 317094 164898 317178 165134
rect 317414 164898 341825 165134
rect 342061 164898 440301 165134
rect 440537 164898 445797 165134
rect 446033 164898 544273 165134
rect 544509 164898 561658 165134
rect 561894 164898 561978 165134
rect 562214 164898 571532 165134
rect 571768 164898 571852 165134
rect 572088 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 9116 147454
rect 9352 147218 9436 147454
rect 9672 147218 31258 147454
rect 31494 147218 31578 147454
rect 31814 147218 58458 147454
rect 58694 147218 58778 147454
rect 59014 147218 85658 147454
rect 85894 147218 85978 147454
rect 86214 147218 112858 147454
rect 113094 147218 113178 147454
rect 113414 147218 140058 147454
rect 140294 147218 140378 147454
rect 140614 147218 167258 147454
rect 167494 147218 167578 147454
rect 167814 147218 194458 147454
rect 194694 147218 194778 147454
rect 195014 147218 221658 147454
rect 221894 147218 221978 147454
rect 222214 147218 248858 147454
rect 249094 147218 249178 147454
rect 249414 147218 276058 147454
rect 276294 147218 276378 147454
rect 276614 147218 303258 147454
rect 303494 147218 303578 147454
rect 303814 147218 330458 147454
rect 330694 147218 330778 147454
rect 331014 147218 357658 147454
rect 357894 147218 357978 147454
rect 358214 147218 384858 147454
rect 385094 147218 385178 147454
rect 385414 147218 412058 147454
rect 412294 147218 412378 147454
rect 412614 147218 439258 147454
rect 439494 147218 439578 147454
rect 439814 147218 466458 147454
rect 466694 147218 466778 147454
rect 467014 147218 493658 147454
rect 493894 147218 493978 147454
rect 494214 147218 520858 147454
rect 521094 147218 521178 147454
rect 521414 147218 548058 147454
rect 548294 147218 548378 147454
rect 548614 147218 570292 147454
rect 570528 147218 570612 147454
rect 570848 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 9116 147134
rect 9352 146898 9436 147134
rect 9672 146898 31258 147134
rect 31494 146898 31578 147134
rect 31814 146898 58458 147134
rect 58694 146898 58778 147134
rect 59014 146898 85658 147134
rect 85894 146898 85978 147134
rect 86214 146898 112858 147134
rect 113094 146898 113178 147134
rect 113414 146898 140058 147134
rect 140294 146898 140378 147134
rect 140614 146898 167258 147134
rect 167494 146898 167578 147134
rect 167814 146898 194458 147134
rect 194694 146898 194778 147134
rect 195014 146898 221658 147134
rect 221894 146898 221978 147134
rect 222214 146898 248858 147134
rect 249094 146898 249178 147134
rect 249414 146898 276058 147134
rect 276294 146898 276378 147134
rect 276614 146898 303258 147134
rect 303494 146898 303578 147134
rect 303814 146898 330458 147134
rect 330694 146898 330778 147134
rect 331014 146898 357658 147134
rect 357894 146898 357978 147134
rect 358214 146898 384858 147134
rect 385094 146898 385178 147134
rect 385414 146898 412058 147134
rect 412294 146898 412378 147134
rect 412614 146898 439258 147134
rect 439494 146898 439578 147134
rect 439814 146898 466458 147134
rect 466694 146898 466778 147134
rect 467014 146898 493658 147134
rect 493894 146898 493978 147134
rect 494214 146898 520858 147134
rect 521094 146898 521178 147134
rect 521414 146898 548058 147134
rect 548294 146898 548378 147134
rect 548614 146898 570292 147134
rect 570528 146898 570612 147134
rect 570848 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 7876 129454
rect 8112 129218 8196 129454
rect 8432 129218 17658 129454
rect 17894 129218 17978 129454
rect 18214 129218 34897 129454
rect 35133 129218 133373 129454
rect 133609 129218 138869 129454
rect 139105 129218 237345 129454
rect 237581 129218 262458 129454
rect 262694 129218 262778 129454
rect 263014 129218 289658 129454
rect 289894 129218 289978 129454
rect 290214 129218 316858 129454
rect 317094 129218 317178 129454
rect 317414 129218 341825 129454
rect 342061 129218 440301 129454
rect 440537 129218 445797 129454
rect 446033 129218 544273 129454
rect 544509 129218 561658 129454
rect 561894 129218 561978 129454
rect 562214 129218 571532 129454
rect 571768 129218 571852 129454
rect 572088 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 7876 129134
rect 8112 128898 8196 129134
rect 8432 128898 17658 129134
rect 17894 128898 17978 129134
rect 18214 128898 34897 129134
rect 35133 128898 133373 129134
rect 133609 128898 138869 129134
rect 139105 128898 237345 129134
rect 237581 128898 262458 129134
rect 262694 128898 262778 129134
rect 263014 128898 289658 129134
rect 289894 128898 289978 129134
rect 290214 128898 316858 129134
rect 317094 128898 317178 129134
rect 317414 128898 341825 129134
rect 342061 128898 440301 129134
rect 440537 128898 445797 129134
rect 446033 128898 544273 129134
rect 544509 128898 561658 129134
rect 561894 128898 561978 129134
rect 562214 128898 571532 129134
rect 571768 128898 571852 129134
rect 572088 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 9116 111454
rect 9352 111218 9436 111454
rect 9672 111218 31258 111454
rect 31494 111218 31578 111454
rect 31814 111218 35617 111454
rect 35853 111218 132653 111454
rect 132889 111218 139589 111454
rect 139825 111218 236625 111454
rect 236861 111218 248858 111454
rect 249094 111218 249178 111454
rect 249414 111218 276058 111454
rect 276294 111218 276378 111454
rect 276614 111218 303258 111454
rect 303494 111218 303578 111454
rect 303814 111218 330458 111454
rect 330694 111218 330778 111454
rect 331014 111218 342545 111454
rect 342781 111218 439581 111454
rect 439817 111218 446517 111454
rect 446753 111218 543553 111454
rect 543789 111218 548058 111454
rect 548294 111218 548378 111454
rect 548614 111218 570292 111454
rect 570528 111218 570612 111454
rect 570848 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 9116 111134
rect 9352 110898 9436 111134
rect 9672 110898 31258 111134
rect 31494 110898 31578 111134
rect 31814 110898 35617 111134
rect 35853 110898 132653 111134
rect 132889 110898 139589 111134
rect 139825 110898 236625 111134
rect 236861 110898 248858 111134
rect 249094 110898 249178 111134
rect 249414 110898 276058 111134
rect 276294 110898 276378 111134
rect 276614 110898 303258 111134
rect 303494 110898 303578 111134
rect 303814 110898 330458 111134
rect 330694 110898 330778 111134
rect 331014 110898 342545 111134
rect 342781 110898 439581 111134
rect 439817 110898 446517 111134
rect 446753 110898 543553 111134
rect 543789 110898 548058 111134
rect 548294 110898 548378 111134
rect 548614 110898 570292 111134
rect 570528 110898 570612 111134
rect 570848 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 7876 93454
rect 8112 93218 8196 93454
rect 8432 93218 17658 93454
rect 17894 93218 17978 93454
rect 18214 93218 34897 93454
rect 35133 93218 133373 93454
rect 133609 93218 138869 93454
rect 139105 93218 237345 93454
rect 237581 93218 262458 93454
rect 262694 93218 262778 93454
rect 263014 93218 289658 93454
rect 289894 93218 289978 93454
rect 290214 93218 316858 93454
rect 317094 93218 317178 93454
rect 317414 93218 341825 93454
rect 342061 93218 440301 93454
rect 440537 93218 445797 93454
rect 446033 93218 544273 93454
rect 544509 93218 561658 93454
rect 561894 93218 561978 93454
rect 562214 93218 571532 93454
rect 571768 93218 571852 93454
rect 572088 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 7876 93134
rect 8112 92898 8196 93134
rect 8432 92898 17658 93134
rect 17894 92898 17978 93134
rect 18214 92898 34897 93134
rect 35133 92898 133373 93134
rect 133609 92898 138869 93134
rect 139105 92898 237345 93134
rect 237581 92898 262458 93134
rect 262694 92898 262778 93134
rect 263014 92898 289658 93134
rect 289894 92898 289978 93134
rect 290214 92898 316858 93134
rect 317094 92898 317178 93134
rect 317414 92898 341825 93134
rect 342061 92898 440301 93134
rect 440537 92898 445797 93134
rect 446033 92898 544273 93134
rect 544509 92898 561658 93134
rect 561894 92898 561978 93134
rect 562214 92898 571532 93134
rect 571768 92898 571852 93134
rect 572088 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 9116 75454
rect 9352 75218 9436 75454
rect 9672 75218 31258 75454
rect 31494 75218 31578 75454
rect 31814 75218 35617 75454
rect 35853 75218 132653 75454
rect 132889 75218 139589 75454
rect 139825 75218 236625 75454
rect 236861 75218 248858 75454
rect 249094 75218 249178 75454
rect 249414 75218 276058 75454
rect 276294 75218 276378 75454
rect 276614 75218 303258 75454
rect 303494 75218 303578 75454
rect 303814 75218 330458 75454
rect 330694 75218 330778 75454
rect 331014 75218 342545 75454
rect 342781 75218 439581 75454
rect 439817 75218 446517 75454
rect 446753 75218 543553 75454
rect 543789 75218 548058 75454
rect 548294 75218 548378 75454
rect 548614 75218 570292 75454
rect 570528 75218 570612 75454
rect 570848 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 9116 75134
rect 9352 74898 9436 75134
rect 9672 74898 31258 75134
rect 31494 74898 31578 75134
rect 31814 74898 35617 75134
rect 35853 74898 132653 75134
rect 132889 74898 139589 75134
rect 139825 74898 236625 75134
rect 236861 74898 248858 75134
rect 249094 74898 249178 75134
rect 249414 74898 276058 75134
rect 276294 74898 276378 75134
rect 276614 74898 303258 75134
rect 303494 74898 303578 75134
rect 303814 74898 330458 75134
rect 330694 74898 330778 75134
rect 331014 74898 342545 75134
rect 342781 74898 439581 75134
rect 439817 74898 446517 75134
rect 446753 74898 543553 75134
rect 543789 74898 548058 75134
rect 548294 74898 548378 75134
rect 548614 74898 570292 75134
rect 570528 74898 570612 75134
rect 570848 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 7876 57454
rect 8112 57218 8196 57454
rect 8432 57218 17658 57454
rect 17894 57218 17978 57454
rect 18214 57218 34897 57454
rect 35133 57218 133373 57454
rect 133609 57218 138869 57454
rect 139105 57218 237345 57454
rect 237581 57218 262458 57454
rect 262694 57218 262778 57454
rect 263014 57218 289658 57454
rect 289894 57218 289978 57454
rect 290214 57218 316858 57454
rect 317094 57218 317178 57454
rect 317414 57218 341825 57454
rect 342061 57218 440301 57454
rect 440537 57218 445797 57454
rect 446033 57218 544273 57454
rect 544509 57218 561658 57454
rect 561894 57218 561978 57454
rect 562214 57218 571532 57454
rect 571768 57218 571852 57454
rect 572088 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 7876 57134
rect 8112 56898 8196 57134
rect 8432 56898 17658 57134
rect 17894 56898 17978 57134
rect 18214 56898 34897 57134
rect 35133 56898 133373 57134
rect 133609 56898 138869 57134
rect 139105 56898 237345 57134
rect 237581 56898 262458 57134
rect 262694 56898 262778 57134
rect 263014 56898 289658 57134
rect 289894 56898 289978 57134
rect 290214 56898 316858 57134
rect 317094 56898 317178 57134
rect 317414 56898 341825 57134
rect 342061 56898 440301 57134
rect 440537 56898 445797 57134
rect 446033 56898 544273 57134
rect 544509 56898 561658 57134
rect 561894 56898 561978 57134
rect 562214 56898 571532 57134
rect 571768 56898 571852 57134
rect 572088 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 9116 39454
rect 9352 39218 9436 39454
rect 9672 39218 31258 39454
rect 31494 39218 31578 39454
rect 31814 39218 58458 39454
rect 58694 39218 58778 39454
rect 59014 39218 85658 39454
rect 85894 39218 85978 39454
rect 86214 39218 112858 39454
rect 113094 39218 113178 39454
rect 113414 39218 140058 39454
rect 140294 39218 140378 39454
rect 140614 39218 167258 39454
rect 167494 39218 167578 39454
rect 167814 39218 194458 39454
rect 194694 39218 194778 39454
rect 195014 39218 221658 39454
rect 221894 39218 221978 39454
rect 222214 39218 248858 39454
rect 249094 39218 249178 39454
rect 249414 39218 276058 39454
rect 276294 39218 276378 39454
rect 276614 39218 303258 39454
rect 303494 39218 303578 39454
rect 303814 39218 330458 39454
rect 330694 39218 330778 39454
rect 331014 39218 357658 39454
rect 357894 39218 357978 39454
rect 358214 39218 384858 39454
rect 385094 39218 385178 39454
rect 385414 39218 412058 39454
rect 412294 39218 412378 39454
rect 412614 39218 439258 39454
rect 439494 39218 439578 39454
rect 439814 39218 466458 39454
rect 466694 39218 466778 39454
rect 467014 39218 493658 39454
rect 493894 39218 493978 39454
rect 494214 39218 520858 39454
rect 521094 39218 521178 39454
rect 521414 39218 548058 39454
rect 548294 39218 548378 39454
rect 548614 39218 570292 39454
rect 570528 39218 570612 39454
rect 570848 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 9116 39134
rect 9352 38898 9436 39134
rect 9672 38898 31258 39134
rect 31494 38898 31578 39134
rect 31814 38898 58458 39134
rect 58694 38898 58778 39134
rect 59014 38898 85658 39134
rect 85894 38898 85978 39134
rect 86214 38898 112858 39134
rect 113094 38898 113178 39134
rect 113414 38898 140058 39134
rect 140294 38898 140378 39134
rect 140614 38898 167258 39134
rect 167494 38898 167578 39134
rect 167814 38898 194458 39134
rect 194694 38898 194778 39134
rect 195014 38898 221658 39134
rect 221894 38898 221978 39134
rect 222214 38898 248858 39134
rect 249094 38898 249178 39134
rect 249414 38898 276058 39134
rect 276294 38898 276378 39134
rect 276614 38898 303258 39134
rect 303494 38898 303578 39134
rect 303814 38898 330458 39134
rect 330694 38898 330778 39134
rect 331014 38898 357658 39134
rect 357894 38898 357978 39134
rect 358214 38898 384858 39134
rect 385094 38898 385178 39134
rect 385414 38898 412058 39134
rect 412294 38898 412378 39134
rect 412614 38898 439258 39134
rect 439494 38898 439578 39134
rect 439814 38898 466458 39134
rect 466694 38898 466778 39134
rect 467014 38898 493658 39134
rect 493894 38898 493978 39134
rect 494214 38898 520858 39134
rect 521094 38898 521178 39134
rect 521414 38898 548058 39134
rect 548294 38898 548378 39134
rect 548614 38898 570292 39134
rect 570528 38898 570612 39134
rect 570848 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 7876 21454
rect 8112 21218 8196 21454
rect 8432 21218 17658 21454
rect 17894 21218 17978 21454
rect 18214 21218 44858 21454
rect 45094 21218 45178 21454
rect 45414 21218 72058 21454
rect 72294 21218 72378 21454
rect 72614 21218 99258 21454
rect 99494 21218 99578 21454
rect 99814 21218 126458 21454
rect 126694 21218 126778 21454
rect 127014 21218 153658 21454
rect 153894 21218 153978 21454
rect 154214 21218 180858 21454
rect 181094 21218 181178 21454
rect 181414 21218 208058 21454
rect 208294 21218 208378 21454
rect 208614 21218 235258 21454
rect 235494 21218 235578 21454
rect 235814 21218 262458 21454
rect 262694 21218 262778 21454
rect 263014 21218 289658 21454
rect 289894 21218 289978 21454
rect 290214 21218 316858 21454
rect 317094 21218 317178 21454
rect 317414 21218 344058 21454
rect 344294 21218 344378 21454
rect 344614 21218 371258 21454
rect 371494 21218 371578 21454
rect 371814 21218 398458 21454
rect 398694 21218 398778 21454
rect 399014 21218 425658 21454
rect 425894 21218 425978 21454
rect 426214 21218 452858 21454
rect 453094 21218 453178 21454
rect 453414 21218 480058 21454
rect 480294 21218 480378 21454
rect 480614 21218 507258 21454
rect 507494 21218 507578 21454
rect 507814 21218 534458 21454
rect 534694 21218 534778 21454
rect 535014 21218 561658 21454
rect 561894 21218 561978 21454
rect 562214 21218 571532 21454
rect 571768 21218 571852 21454
rect 572088 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 7876 21134
rect 8112 20898 8196 21134
rect 8432 20898 17658 21134
rect 17894 20898 17978 21134
rect 18214 20898 44858 21134
rect 45094 20898 45178 21134
rect 45414 20898 72058 21134
rect 72294 20898 72378 21134
rect 72614 20898 99258 21134
rect 99494 20898 99578 21134
rect 99814 20898 126458 21134
rect 126694 20898 126778 21134
rect 127014 20898 153658 21134
rect 153894 20898 153978 21134
rect 154214 20898 180858 21134
rect 181094 20898 181178 21134
rect 181414 20898 208058 21134
rect 208294 20898 208378 21134
rect 208614 20898 235258 21134
rect 235494 20898 235578 21134
rect 235814 20898 262458 21134
rect 262694 20898 262778 21134
rect 263014 20898 289658 21134
rect 289894 20898 289978 21134
rect 290214 20898 316858 21134
rect 317094 20898 317178 21134
rect 317414 20898 344058 21134
rect 344294 20898 344378 21134
rect 344614 20898 371258 21134
rect 371494 20898 371578 21134
rect 371814 20898 398458 21134
rect 398694 20898 398778 21134
rect 399014 20898 425658 21134
rect 425894 20898 425978 21134
rect 426214 20898 452858 21134
rect 453094 20898 453178 21134
rect 453414 20898 480058 21134
rect 480294 20898 480378 21134
rect 480614 20898 507258 21134
rect 507494 20898 507578 21134
rect 507814 20898 534458 21134
rect 534694 20898 534778 21134
rect 535014 20898 561658 21134
rect 561894 20898 561978 21134
rect 562214 20898 571532 21134
rect 571768 20898 571852 21134
rect 572088 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use user_proj_example  mprj
timestamp 0
transform 1 0 4000 0 1 4000
box 0 0 571964 694008
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 2000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 700008 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 700008 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 700008 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 700008 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 700008 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 700008 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 700008 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 700008 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 700008 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 700008 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 700008 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 700008 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 700008 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 700008 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 700008 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 700008 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 700008 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 2000 8 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 700008 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 700008 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 700008 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 700008 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 700008 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 700008 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 700008 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 700008 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 700008 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 700008 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 700008 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 700008 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 700008 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 700008 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 700008 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 700008 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 2000 8 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 700008 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 700008 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 700008 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 700008 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 700008 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 700008 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 700008 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 700008 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 700008 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 700008 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 700008 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 700008 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 700008 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 700008 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 700008 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 700008 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 2000 8 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 700008 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 700008 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 700008 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 700008 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 700008 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 700008 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 700008 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 700008 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 700008 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 700008 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 700008 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 700008 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 700008 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 700008 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 700008 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 700008 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 700008 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 700008 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 700008 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 700008 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 700008 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 700008 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 700008 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 700008 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 700008 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 700008 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 700008 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 700008 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 700008 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 700008 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 700008 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 700008 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 700008 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 700008 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 700008 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 700008 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 700008 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 700008 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 700008 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 700008 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 700008 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 700008 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 700008 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 700008 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 700008 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 700008 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 700008 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 700008 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 2000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 700008 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 700008 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 700008 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 700008 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 700008 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 700008 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 700008 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 700008 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 700008 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 700008 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 700008 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 700008 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 700008 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 700008 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 700008 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 700008 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 700008 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 700008 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 700008 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 700008 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 700008 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 700008 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 700008 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 700008 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 700008 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 700008 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 700008 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 700008 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 700008 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 700008 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 700008 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 700008 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
